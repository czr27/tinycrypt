--
-- SKINNY-AEAD Reference Hardware Implementation
-- 
-- Copyright 2019:
--     Amir Moradi & Pascal Sasdrich for the SKINNY Team
--     https://sites.google.com/site/skinnycipher/
-- 
-- This program is free software; you can redistribute it and/or
-- modify it under the terms of the GNU General Public License as
-- published by the Free Software Foundation; either version 2 of the
-- License, or (at your option) any later version.
-- 
-- This program is distributed in the hope that it will be useful, but
-- WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE. See the GNU
-- General Public License for more details.
-- 

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE IEEE.std_logic_textio.all;
USE ieee.numeric_std.ALL;
USE ieee.math_real.ALL; 

ENTITY SKINNY_tk3_AEAD_encdec_M1_Test_Part1 IS
END SKINNY_tk3_AEAD_encdec_M1_Test_Part1;
 
ARCHITECTURE behavior OF SKINNY_tk3_AEAD_encdec_M1_Test_Part1 IS 
 
	constant	nl		 : integer := 0; -- 128-bit nonce
	constant	tl		 : integer := 0; -- 128-bit tag     -> M1
 
 
   COMPONENT SKINNY_tk3_AEAD
	Generic (
		nl				 : integer;  -- 0: 128-bit nonce, 1: 96-bit nonce
		tl				 : integer); -- 0: 128-bit tag,   1: 64-bit tag
	Port (  
		clk          : in  STD_LOGIC;
		rst      	 : in  STD_LOGIC;
		a_data       : in  STD_LOGIC;
		enc          : in  STD_LOGIC;
		dec          : in  STD_LOGIC;
		gen_tag      : in  std_logic;
		Input1       : in  STD_LOGIC_VECTOR (127       downto 0);  -- Message or Associated Data (share 1)
		Input2       : in  STD_LOGIC_VECTOR (127       downto 0);  -- Message or Associated Data (share 2)
		N            : in  STD_LOGIC_VECTOR (127-nl*32 downto 0);
		K1           : in  STD_LOGIC_VECTOR (127       downto 0); -- Key (share 1)
		K2           : in  STD_LOGIC_VECTOR (127       downto 0); -- Key (share 2)
		Block_Size	 : in  STD_LOGIC_VECTOR (  3       downto 0); -- Size of the given block as Input (in BYTES) - 1
		Output1      : out STD_LOGIC_VECTOR (127       downto 0); -- Ciphertext (share 1)
		Output2      : out STD_LOGIC_VECTOR (127       downto 0); -- Ciphertext (share 2) 
		Tag1			 : out STD_LOGIC_VECTOR (127-tl*64 downto 0); -- Tag (share 1)
		Tag2			 : out STD_LOGIC_VECTOR (127-tl*64 downto 0); -- Tag (share 2)
		done         : out STD_LOGIC);
	END COMPONENT;
    

   --Inputs
   signal clk 			: std_logic := '0';
   signal rst 			: std_logic := '0';
   signal a_data 		: std_logic := '0';
   signal enc 			: std_logic := '0';
   signal dec 			: std_logic := '0';
   signal gen_tag 	: std_logic := '0';
   signal Input1 		: std_logic_vector(127       downto 0) := (others => '0');
   signal Input2 		: std_logic_vector(127       downto 0) := (others => '0');
   signal N 			: std_logic_vector(127-nl*32 downto 0) := (others => '0');
   signal K1 			: std_logic_vector(127       downto 0) := (others => '0');
   signal K2 			: std_logic_vector(127       downto 0) := (others => '0');
   signal Block_Size : std_logic_vector(  3       downto 0) := (others => '0');

 	--Outputs
   signal Output1		: std_logic_vector(127 downto 0);
   signal Output2		: std_logic_vector(127 downto 0);
   signal Tag1		   : std_logic_vector(127-tl*64 downto 0);
   signal Tag2		   : std_logic_vector(127-tl*64 downto 0);
   signal done 		: std_logic;

   signal Input 		: std_logic_vector(127 downto 0) := (others => '0');
   signal K 			: std_logic_vector(127 downto 0) := (others => '0');
   signal Output		: std_logic_vector(127 downto 0);
   signal Tag		   : std_logic_vector(127-tl*64 downto 0);

	signal Mask1		: std_logic_vector(127 downto 0);
	signal Mask2		: std_logic_vector(127 downto 0);
	

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
 	type INT_ARRAY  is array (integer range <>) of integer range 0 to 255;
	type REAL_ARRAY is array (integer range <>) of real;
	type BYTE_ARRAY is array (integer range <>) of std_logic_vector(7 downto 0);

	signal r: INT_ARRAY (31 downto 0);
	signal m: BYTE_ARRAY(31 downto 0);

BEGIN
 
  	maskgen: process
		 variable seed1, seed2: positive;        -- seed values for random generator
		 variable rand: REAL_ARRAY(31 downto 0); -- random real-number value in range 0 to 1.0  
		 variable range_of_rand : real := 256.0; -- the range of random values created will be 0 to +255.
	begin
		 
		FOR i in 0 to 31 loop
			uniform(seed1, seed2, rand(i));   -- generate random number
			r(i) <= integer(TRUNC(rand(i)*range_of_rand));  -- rescale to 0...255, convert integer part 
			m(i) <= std_logic_vector(to_unsigned(r(i), m(i)'length));
		end loop;
		
		wait for clk_period;
	end process;  

	---------
	
	maskassign: FOR i in 0 to 15 GENERATE
		Mask1(i*8+7 downto i*8)	<= m(i);
		Mask2(i*8+7 downto i*8)	<= m(16+i);
	END GENERATE;

	---------
 
   uut: SKINNY_tk3_AEAD 
	GENERIC MAP (
		nl		=> nl,
		tl		=> tl)
	PORT MAP (
		clk 			=> clk,
		rst 			=> rst,
		a_data 		=> a_data,
		enc 			=> enc,
		dec			=> dec,
		gen_tag 		=> gen_tag,
		Input1 		=> Input1,
		Input2 		=> Input2,
		N 				=> N,
		K1				=> K1,
		K2				=> K2,
		Block_Size 	=> Block_Size,
		Output1 		=> Output1,
		Output2 		=> Output2,
		Tag1			=> Tag1,
		Tag2			=> Tag2,
		done 			=> done);

	Input1	<= Input XOR Mask1;
	Input2	<= Mask1;

	K1			<= K XOR Mask2;
	K2			<= Mask2;

	Output	<= Output1 XOR Output2;
	Tag		<= Tag1 XOR Tag2;


   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      --------- test no. 1 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"99CE68EF7B52AAD0E11C6E2FC722426D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 2 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4720E8EA3682D9E9DC5C83563705F8F4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 3 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"66082EC45370954D65EB5A06B35D992B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 4 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C29FDF3EEB81A8314859230542FC45B4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 5 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CA192E010E95F8A309DE331261B83887") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 6 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DE8A628D49B00A8F70C1C87A89CE622D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 7 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EAF7736E366F6D8BC2E9CD7FDA8B8A7F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 8 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D77102862CABCDEB212F1F88360357EF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 9 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FA83E300D6C9FC7B24ABF86AD7F2F221") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 10 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CBF0269A295608E3801F3FFFD1571161") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 11 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"386C476D3BDA8CBD205B50AFF2D12E6E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 12 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0370ACA4142DFBFBCCF3FED1CAF17CDA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 13 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F8A1E33C1B60E68C1777B8376FDCA936") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 14 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"72CD0A85F19AF6F6D1FDB4ACFF66FCA9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 15 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"43175F8DF12BB951396DAB712ECD582F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 16 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C6CB80856D50604735D970FA5488FF23") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 17 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"764ADBD8C65326C00DFF319C5D23B7FD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 18 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C84CE30DF583E4C0F582560E64643C17") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 19 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F7E217673E83BAEB5325E5E739C612AA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 20 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6F956F4D1E93E1192F3BF339E248617A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 21 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"13A38E78FA2D2AB63249E4AEFC3BB4CD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 22 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1343DEA3E2891FB20352A64D7440729F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 23 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C0BA4F75568F44C029101E5D96CCBA10") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 24 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"06AF4F6F56C0A4A3818FA83F97508D92") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 25 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"80B61783EBB692B86255879BB04BB304") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 26 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2BCDC384E3CFD5C3D7198F949C471574") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 27 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"32A9DD75E2BA0E137383D3EEE2A07E34") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 28 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"877927B4EC6E76D543E6AAB2BE235907") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 29 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4907500E302AE30B4547C47E9D046A45") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 30 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F3FC1A3B7A89B1AD26BEFD26C8E5B14E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 31 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5047617083F872D7F75DDAFDA8D1C24B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 32 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"08F611836F47F00286D7EB25DC1BB620") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 33 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"363BA410E56D196796761F338410F6AF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 34 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"85") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C6E991B30CC1479902E0E9736CA436F6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"85";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C6E991B30CC1479902E0E9736CA436F6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 35 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"85") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"180711B6411134A03FA0040A9C838C6F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"85";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"180711B6411134A03FA0040A9C838C6F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 36 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"85") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"392FD79824E378048617DD5A18DBEDB0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"85";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"392FD79824E378048617DD5A18DBEDB0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 37 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"85") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9DB826629C124578ABA5A459E97A312F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"85";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9DB826629C124578ABA5A459E97A312F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 38 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"85") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"953ED75D790615EAEA22B44ECA3E4C1C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"85";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"953ED75D790615EAEA22B44ECA3E4C1C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 39 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"85") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"81AD9BD13E23E7C6933D4F26224816B6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"85";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"81AD9BD13E23E7C6933D4F26224816B6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 40 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"85") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B5D08A3241FC80C221154A23710DFEE4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"85";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B5D08A3241FC80C221154A23710DFEE4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 41 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"85") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8856FBDA5B3820A2C2D398D49D852374") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"85";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8856FBDA5B3820A2C2D398D49D852374") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 42 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"85") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A5A41A5CA15A1132C7577F367C7486BA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"85";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A5A41A5CA15A1132C7577F367C7486BA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 43 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"85") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"94D7DFC65EC5E5AA63E3B8A37AD165FA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"85";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"94D7DFC65EC5E5AA63E3B8A37AD165FA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 44 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"85") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"674BBE314C4961F4C3A7D7F359575AF5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"85";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"674BBE314C4961F4C3A7D7F359575AF5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 45 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"85") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5C5755F863BE16B22F0F798D61770841") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"85";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5C5755F863BE16B22F0F798D61770841") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 46 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"85") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A7861A606CF30BC5F48B3F6BC45ADDAD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"85";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A7861A606CF30BC5F48B3F6BC45ADDAD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 47 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"85") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2DEAF3D986091BBF320133F054E08832") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"85";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2DEAF3D986091BBF320133F054E08832") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 48 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"85") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1C30A6D186B85418DA912C2D854B2CB4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"85";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1C30A6D186B85418DA912C2D854B2CB4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 49 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"85") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"99EC79D91AC38D0ED625F7A6FF0E8BB8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"85";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"99EC79D91AC38D0ED625F7A6FF0E8BB8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 50 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"85") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"296D2284B1C0CB89EE03B6C0F6A5C366") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"85";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"296D2284B1C0CB89EE03B6C0F6A5C366") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 51 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"85") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"976B1A5182100989167ED152CFE2488C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"85";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"976B1A5182100989167ED152CFE2488C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 52 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"85") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A8C5EE3B491057A2B0D962BB92406631") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"85";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A8C5EE3B491057A2B0D962BB92406631") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 53 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"85") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"30B2961169000C50CCC7746549CE15E1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"85";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"30B2961169000C50CCC7746549CE15E1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 54 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"85") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4C8477248DBEC7FFD1B563F257BDC056") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"85";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4C8477248DBEC7FFD1B563F257BDC056") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 55 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"85") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4C6427FF951AF2FBE0AE2111DFC60604") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"85";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4C6427FF951AF2FBE0AE2111DFC60604") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 56 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"85") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9F9DB629211CA989CAEC99013D4ACE8B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"85";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9F9DB629211CA989CAEC99013D4ACE8B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 57 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"85") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5988B633215349EA62732F633CD6F909") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"85";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5988B633215349EA62732F633CD6F909") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 58 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"85") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DF91EEDF9C257FF181A900C71BCDC79F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"85";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DF91EEDF9C257FF181A900C71BCDC79F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 59 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"85") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"74EA3AD8945C388A34E508C837C161EF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"85";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"74EA3AD8945C388A34E508C837C161EF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 60 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"85") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6D8E24299529E35A907F54B249260AAF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"85";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6D8E24299529E35A907F54B249260AAF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 61 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"85") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D85EDEE89BFD9B9CA01A2DEE15A52D9C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"85";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D85EDEE89BFD9B9CA01A2DEE15A52D9C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 62 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"85") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1620A95247B90E42A6BB432236821EDE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"85";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1620A95247B90E42A6BB432236821EDE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 63 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"85") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"ACDBE3670D1A5CE4C5427A7A6363C5D5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"85";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"ACDBE3670D1A5CE4C5427A7A6363C5D5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 64 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"85") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0F60982CF46B9F9E14A15DA10357B6D0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"85";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0F60982CF46B9F9E14A15DA10357B6D0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 65 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"85") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"57D1E8DF18D41D4B652B6C79779DC2BB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"85";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"57D1E8DF18D41D4B652B6C79779DC2BB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 66 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"85") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"691C5D4C92FEF42E758A986F2F968234") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"85";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"691C5D4C92FEF42E758A986F2F968234") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 67 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"85BB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CE4030AA00B908B523BF711D27013807") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"85BB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CE4030AA00B908B523BF711D27013807") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 68 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"85BB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"10AEB0AF4D697B8C1EFF9C64D726829E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"85BB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"10AEB0AF4D697B8C1EFF9C64D726829E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 69 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"85BB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"31867681289B3728A7484534537EE341") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"85BB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"31867681289B3728A7484534537EE341") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 70 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"85BB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9511877B906A0A548AFA3C37A2DF3FDE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"85BB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9511877B906A0A548AFA3C37A2DF3FDE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 71 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"85BB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9D977644757E5AC6CB7D2C20819B42ED") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"85BB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9D977644757E5AC6CB7D2C20819B42ED") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 72 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"85BB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"89043AC8325BA8EAB262D74869ED1847") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"85BB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"89043AC8325BA8EAB262D74869ED1847") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 73 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"85BB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BD792B2B4D84CFEE004AD24D3AA8F015") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"85BB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BD792B2B4D84CFEE004AD24D3AA8F015") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 74 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"85BB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"80FF5AC357406F8EE38C00BAD6202D85") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"85BB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"80FF5AC357406F8EE38C00BAD6202D85") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 75 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"85BB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AD0DBB45AD225E1EE608E75837D1884B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"85BB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AD0DBB45AD225E1EE608E75837D1884B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 76 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"85BB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9C7E7EDF52BDAA8642BC20CD31746B0B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"85BB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9C7E7EDF52BDAA8642BC20CD31746B0B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 77 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"85BB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6FE21F2840312ED8E2F84F9D12F25404") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"85BB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6FE21F2840312ED8E2F84F9D12F25404") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 78 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"85BB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"54FEF4E16FC6599E0E50E1E32AD206B0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"85BB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"54FEF4E16FC6599E0E50E1E32AD206B0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 79 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"85BB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AF2FBB79608B44E9D5D4A7058FFFD35C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"85BB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AF2FBB79608B44E9D5D4A7058FFFD35C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 80 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"85BB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"254352C08A715493135EAB9E1F4586C3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"85BB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"254352C08A715493135EAB9E1F4586C3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 81 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"85BB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"149907C88AC01B34FBCEB443CEEE2245") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"85BB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"149907C88AC01B34FBCEB443CEEE2245") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 82 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"85BB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9145D8C016BBC222F77A6FC8B4AB8549") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"85BB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9145D8C016BBC222F77A6FC8B4AB8549") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 83 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"85BB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"21C4839DBDB884A5CF5C2EAEBD00CD97") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"85BB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"21C4839DBDB884A5CF5C2EAEBD00CD97") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 84 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"85BB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9FC2BB488E6846A53721493C8447467D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"85BB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9FC2BB488E6846A53721493C8447467D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 85 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"85BB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A06C4F224568188E9186FAD5D9E568C0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"85BB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A06C4F224568188E9186FAD5D9E568C0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 86 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"85BB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"381B37086578437CED98EC0B026B1B10") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"85BB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"381B37086578437CED98EC0B026B1B10") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 87 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"85BB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"442DD63D81C688D3F0EAFB9C1C18CEA7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"85BB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"442DD63D81C688D3F0EAFB9C1C18CEA7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 88 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"85BB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"44CD86E69962BDD7C1F1B97F946308F5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"85BB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"44CD86E69962BDD7C1F1B97F946308F5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 89 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"85BB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"973417302D64E6A5EBB3016F76EFC07A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"85BB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"973417302D64E6A5EBB3016F76EFC07A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 90 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"85BB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5121172A2D2B06C6432CB70D7773F7F8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"85BB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5121172A2D2B06C6432CB70D7773F7F8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 91 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"85BB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D7384FC6905D30DDA0F698A95068C96E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"85BB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D7384FC6905D30DDA0F698A95068C96E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 92 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"85BB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7C439BC1982477A615BA90A67C646F1E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"85BB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7C439BC1982477A615BA90A67C646F1E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 93 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"85BB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"652785309951AC76B120CCDC0283045E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"85BB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"652785309951AC76B120CCDC0283045E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 94 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"85BB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D0F77FF19785D4B08145B5805E00236D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"85BB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D0F77FF19785D4B08145B5805E00236D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 95 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"85BB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1E89084B4BC1416E87E4DB4C7D27102F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"85BB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1E89084B4BC1416E87E4DB4C7D27102F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 96 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"85BB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A472427E016213C8E41DE21428C6CB24") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"85BB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A472427E016213C8E41DE21428C6CB24") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 97 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"85BB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"07C93935F813D0B235FEC5CF48F2B821") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"85BB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"07C93935F813D0B235FEC5CF48F2B821") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 98 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"85BB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5F7849C614AC52674474F4173C38CC4A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"85BB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5F7849C614AC52674474F4173C38CC4A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 99 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"85BB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"61B5FC559E86BB0254D5000164338CC5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"85BB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"61B5FC559E86BB0254D5000164338CC5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 100 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"85BBEA") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"90928187998C34F5D5FB5A50B8FCE96D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"85BBEA";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"90928187998C34F5D5FB5A50B8FCE96D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 101 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"85BBEA") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4E7C0182D45C47CCE8BBB72948DB53F4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"85BBEA";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4E7C0182D45C47CCE8BBB72948DB53F4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 102 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"85BBEA") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6F54C7ACB1AE0B68510C6E79CC83322B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"85BBEA";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6F54C7ACB1AE0B68510C6E79CC83322B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 103 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"85BBEA") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CBC33656095F36147CBE177A3D22EEB4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"85BBEA";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CBC33656095F36147CBE177A3D22EEB4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 104 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"85BBEA") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C345C769EC4B66863D39076D1E669387") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"85BBEA";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C345C769EC4B66863D39076D1E669387") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 105 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"85BBEA") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D7D68BE5AB6E94AA4426FC05F610C92D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"85BBEA";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D7D68BE5AB6E94AA4426FC05F610C92D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 106 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"85BBEA") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E3AB9A06D4B1F3AEF60EF900A555217F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"85BBEA";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E3AB9A06D4B1F3AEF60EF900A555217F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 107 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"85BBEA") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DE2DEBEECE7553CE15C82BF749DDFCEF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"85BBEA";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DE2DEBEECE7553CE15C82BF749DDFCEF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 108 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"85BBEA") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F3DF0A683417625E104CCC15A82C5921") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"85BBEA";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F3DF0A683417625E104CCC15A82C5921") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 109 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"85BBEA") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C2ACCFF2CB8896C6B4F80B80AE89BA61") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"85BBEA";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C2ACCFF2CB8896C6B4F80B80AE89BA61") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 110 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"85BBEA") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3130AE05D904129814BC64D08D0F856E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"85BBEA";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3130AE05D904129814BC64D08D0F856E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 111 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"85BBEA") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0A2C45CCF6F365DEF814CAAEB52FD7DA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"85BBEA";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0A2C45CCF6F365DEF814CAAEB52FD7DA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 112 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"85BBEA") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F1FD0A54F9BE78A923908C4810020236") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"85BBEA";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F1FD0A54F9BE78A923908C4810020236") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 113 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"85BBEA") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7B91E3ED134468D3E51A80D380B857A9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"85BBEA";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7B91E3ED134468D3E51A80D380B857A9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 114 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"85BBEA") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4A4BB6E513F527740D8A9F0E5113F32F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"85BBEA";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4A4BB6E513F527740D8A9F0E5113F32F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 115 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"85BBEA") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CF9769ED8F8EFE62013E44852B565423") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"85BBEA";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CF9769ED8F8EFE62013E44852B565423") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 116 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"85BBEA") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7F1632B0248DB8E5391805E322FD1CFD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"85BBEA";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7F1632B0248DB8E5391805E322FD1CFD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 117 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"85BBEA") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C1100A65175D7AE5C16562711BBA9717") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"85BBEA";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C1100A65175D7AE5C16562711BBA9717") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 118 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"85BBEA") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FEBEFE0FDC5D24CE67C2D1984618B9AA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"85BBEA";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FEBEFE0FDC5D24CE67C2D1984618B9AA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 119 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"85BBEA") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"66C98625FC4D7F3C1BDCC7469D96CA7A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"85BBEA";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"66C98625FC4D7F3C1BDCC7469D96CA7A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 120 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"85BBEA") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1AFF671018F3B49306AED0D183E51FCD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"85BBEA";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1AFF671018F3B49306AED0D183E51FCD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 121 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"85BBEA") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1A1F37CB0057819737B592320B9ED99F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"85BBEA";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1A1F37CB0057819737B592320B9ED99F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 122 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"85BBEA") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C9E6A61DB451DAE51DF72A22E9121110") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"85BBEA";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C9E6A61DB451DAE51DF72A22E9121110") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 123 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"85BBEA") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0FF3A607B41E3A86B5689C40E88E2692") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"85BBEA";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0FF3A607B41E3A86B5689C40E88E2692") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 124 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"85BBEA") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"89EAFEEB09680C9D56B2B3E4CF951804") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"85BBEA";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"89EAFEEB09680C9D56B2B3E4CF951804") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 125 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"85BBEA") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"22912AEC01114BE6E3FEBBEBE399BE74") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"85BBEA";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"22912AEC01114BE6E3FEBBEBE399BE74") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 126 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"85BBEA") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3BF5341D006490364764E7919D7ED534") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"85BBEA";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3BF5341D006490364764E7919D7ED534") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 127 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"85BBEA") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8E25CEDC0EB0E8F077019ECDC1FDF207") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"85BBEA";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8E25CEDC0EB0E8F077019ECDC1FDF207") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 128 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"85BBEA") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"405BB966D2F47D2E71A0F001E2DAC145") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"85BBEA";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"405BB966D2F47D2E71A0F001E2DAC145") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 129 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"85BBEA") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FAA0F35398572F881259C959B73B1A4E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"85BBEA";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FAA0F35398572F881259C959B73B1A4E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 130 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"85BBEA") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"591B88186126ECF2C3BAEE82D70F694B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"85BBEA";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"591B88186126ECF2C3BAEE82D70F694B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 131 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"85BBEA") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"01AAF8EB8D996E27B230DF5AA3C51D20") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"85BBEA";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"01AAF8EB8D996E27B230DF5AA3C51D20") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 132 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"85BBEA") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3F674D7807B38742A2912B4CFBCE5DAF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"85BBEA";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3F674D7807B38742A2912B4CFBCE5DAF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 133 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"85BBEAE2") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C4F64ABC86580C2E4CD19A2E9655165F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"85BBEAE2";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C4F64ABC86580C2E4CD19A2E9655165F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 134 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"85BBEAE2") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1A18CAB9CB887F17719177576672ACC6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"85BBEAE2";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1A18CAB9CB887F17719177576672ACC6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 135 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"85BBEAE2") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3B300C97AE7A33B3C826AE07E22ACD19") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"85BBEAE2";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3B300C97AE7A33B3C826AE07E22ACD19") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 136 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"85BBEAE2") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9FA7FD6D168B0ECFE594D704138B1186") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"85BBEAE2";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9FA7FD6D168B0ECFE594D704138B1186") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 137 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"85BBEAE2") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"97210C52F39F5E5DA413C71330CF6CB5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"85BBEAE2";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"97210C52F39F5E5DA413C71330CF6CB5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 138 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"85BBEAE2") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"83B240DEB4BAAC71DD0C3C7BD8B9361F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"85BBEAE2";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"83B240DEB4BAAC71DD0C3C7BD8B9361F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 139 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"85BBEAE2") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B7CF513DCB65CB756F24397E8BFCDE4D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"85BBEAE2";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B7CF513DCB65CB756F24397E8BFCDE4D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 140 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"85BBEAE2") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8A4920D5D1A16B158CE2EB89677403DD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"85BBEAE2";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8A4920D5D1A16B158CE2EB89677403DD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 141 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"85BBEAE2") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A7BBC1532BC35A8589660C6B8685A613") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"85BBEAE2";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A7BBC1532BC35A8589660C6B8685A613") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 142 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"85BBEAE2") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"96C804C9D45CAE1D2DD2CBFE80204553") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"85BBEAE2";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"96C804C9D45CAE1D2DD2CBFE80204553") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 143 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"85BBEAE2") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6554653EC6D02A438D96A4AEA3A67A5C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"85BBEAE2";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6554653EC6D02A438D96A4AEA3A67A5C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 144 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"85BBEAE2") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5E488EF7E9275D05613E0AD09B8628E8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"85BBEAE2";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5E488EF7E9275D05613E0AD09B8628E8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 145 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"85BBEAE2") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A599C16FE66A4072BABA4C363EABFD04") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"85BBEAE2";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A599C16FE66A4072BABA4C363EABFD04") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 146 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"85BBEAE2") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2FF528D60C9050087C3040ADAE11A89B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"85BBEAE2";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2FF528D60C9050087C3040ADAE11A89B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 147 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"85BBEAE2") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1E2F7DDE0C211FAF94A05F707FBA0C1D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"85BBEAE2";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1E2F7DDE0C211FAF94A05F707FBA0C1D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 148 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"85BBEAE2") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9BF3A2D6905AC6B9981484FB05FFAB11") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"85BBEAE2";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9BF3A2D6905AC6B9981484FB05FFAB11") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 149 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"85BBEAE2") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2B72F98B3B59803EA032C59D0C54E3CF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"85BBEAE2";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2B72F98B3B59803EA032C59D0C54E3CF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 150 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"85BBEAE2") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9574C15E0889423E584FA20F35136825") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"85BBEAE2";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9574C15E0889423E584FA20F35136825") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 151 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"85BBEAE2") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AADA3534C3891C15FEE811E668B14698") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"85BBEAE2";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AADA3534C3891C15FEE811E668B14698") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 152 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"85BBEAE2") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"32AD4D1EE39947E782F60738B33F3548") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"85BBEAE2";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"32AD4D1EE39947E782F60738B33F3548") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 153 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"85BBEAE2") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4E9BAC2B07278C489F8410AFAD4CE0FF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"85BBEAE2";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4E9BAC2B07278C489F8410AFAD4CE0FF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 154 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"85BBEAE2") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4E7BFCF01F83B94CAE9F524C253726AD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"85BBEAE2";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4E7BFCF01F83B94CAE9F524C253726AD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 155 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"85BBEAE2") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9D826D26AB85E23E84DDEA5CC7BBEE22") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"85BBEAE2";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9D826D26AB85E23E84DDEA5CC7BBEE22") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 156 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"85BBEAE2") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5B976D3CABCA025D2C425C3EC627D9A0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"85BBEAE2";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5B976D3CABCA025D2C425C3EC627D9A0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 157 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"85BBEAE2") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DD8E35D016BC3446CF98739AE13CE736") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"85BBEAE2";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DD8E35D016BC3446CF98739AE13CE736") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 158 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"85BBEAE2") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"76F5E1D71EC5733D7AD47B95CD304146") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"85BBEAE2";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"76F5E1D71EC5733D7AD47B95CD304146") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 159 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"85BBEAE2") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6F91FF261FB0A8EDDE4E27EFB3D72A06") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"85BBEAE2";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6F91FF261FB0A8EDDE4E27EFB3D72A06") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 160 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"85BBEAE2") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DA4105E71164D02BEE2B5EB3EF540D35") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"85BBEAE2";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DA4105E71164D02BEE2B5EB3EF540D35") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 161 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"85BBEAE2") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"143F725DCD2045F5E88A307FCC733E77") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"85BBEAE2";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"143F725DCD2045F5E88A307FCC733E77") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 162 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"85BBEAE2") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AEC43868878317538B7309279992E57C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"85BBEAE2";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AEC43868878317538B7309279992E57C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 163 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"85BBEAE2") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0D7F43237EF2D4295A902EFCF9A69679") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"85BBEAE2";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0D7F43237EF2D4295A902EFCF9A69679") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 164 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"85BBEAE2") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"55CE33D0924D56FC2B1A1F248D6CE212") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"85BBEAE2";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"55CE33D0924D56FC2B1A1F248D6CE212") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 165 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"85BBEAE2") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6B0386431867BF993BBBEB32D567A29D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"85BBEAE2";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6B0386431867BF993BBBEB32D567A29D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 166 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"85BBEAE208") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0F697EFF63AC2A88CD6A13AC069A117D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"85BBEAE208";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0F697EFF63AC2A88CD6A13AC069A117D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 167 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"85BBEAE208") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D187FEFA2E7C59B1F02AFED5F6BDABE4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"85BBEAE208";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D187FEFA2E7C59B1F02AFED5F6BDABE4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 168 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"85BBEAE208") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F0AF38D44B8E1515499D278572E5CA3B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"85BBEAE208";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F0AF38D44B8E1515499D278572E5CA3B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 169 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"85BBEAE208") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5438C92EF37F2869642F5E86834416A4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"85BBEAE208";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5438C92EF37F2869642F5E86834416A4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 170 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"85BBEAE208") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5CBE3811166B78FB25A84E91A0006B97") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"85BBEAE208";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5CBE3811166B78FB25A84E91A0006B97") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 171 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"85BBEAE208") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"482D749D514E8AD75CB7B5F94876313D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"85BBEAE208";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"482D749D514E8AD75CB7B5F94876313D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 172 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"85BBEAE208") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7C50657E2E91EDD3EE9FB0FC1B33D96F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"85BBEAE208";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7C50657E2E91EDD3EE9FB0FC1B33D96F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 173 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"85BBEAE208") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"41D6149634554DB30D59620BF7BB04FF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"85BBEAE208";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"41D6149634554DB30D59620BF7BB04FF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 174 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"85BBEAE208") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6C24F510CE377C2308DD85E9164AA131") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"85BBEAE208";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6C24F510CE377C2308DD85E9164AA131") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 175 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"85BBEAE208") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5D57308A31A888BBAC69427C10EF4271") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"85BBEAE208";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5D57308A31A888BBAC69427C10EF4271") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 176 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"85BBEAE208") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AECB517D23240CE50C2D2D2C33697D7E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"85BBEAE208";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AECB517D23240CE50C2D2D2C33697D7E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 177 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"85BBEAE208") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"95D7BAB40CD37BA3E08583520B492FCA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"85BBEAE208";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"95D7BAB40CD37BA3E08583520B492FCA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 178 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"85BBEAE208") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6E06F52C039E66D43B01C5B4AE64FA26") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"85BBEAE208";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6E06F52C039E66D43B01C5B4AE64FA26") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 179 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"85BBEAE208") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E46A1C95E96476AEFD8BC92F3EDEAFB9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"85BBEAE208";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E46A1C95E96476AEFD8BC92F3EDEAFB9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 180 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"85BBEAE208") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D5B0499DE9D53909151BD6F2EF750B3F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"85BBEAE208";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D5B0499DE9D53909151BD6F2EF750B3F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 181 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"85BBEAE208") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"506C969575AEE01F19AF0D799530AC33") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"85BBEAE208";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"506C969575AEE01F19AF0D799530AC33") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 182 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"85BBEAE208") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E0EDCDC8DEADA69821894C1F9C9BE4ED") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"85BBEAE208";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E0EDCDC8DEADA69821894C1F9C9BE4ED") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 183 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"85BBEAE208") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5EEBF51DED7D6498D9F42B8DA5DC6F07") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"85BBEAE208";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5EEBF51DED7D6498D9F42B8DA5DC6F07") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 184 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"85BBEAE208") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"61450177267D3AB37F539864F87E41BA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"85BBEAE208";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"61450177267D3AB37F539864F87E41BA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 185 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"85BBEAE208") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F932795D066D6141034D8EBA23F0326A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"85BBEAE208";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F932795D066D6141034D8EBA23F0326A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 186 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"85BBEAE208") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"85049868E2D3AAEE1E3F992D3D83E7DD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"85BBEAE208";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"85049868E2D3AAEE1E3F992D3D83E7DD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 187 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"85BBEAE208") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"85E4C8B3FA779FEA2F24DBCEB5F8218F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"85BBEAE208";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"85E4C8B3FA779FEA2F24DBCEB5F8218F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 188 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"85BBEAE208") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"561D59654E71C498056663DE5774E900") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"85BBEAE208";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"561D59654E71C498056663DE5774E900") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 189 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"85BBEAE208") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9008597F4E3E24FBADF9D5BC56E8DE82") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"85BBEAE208";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9008597F4E3E24FBADF9D5BC56E8DE82") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 190 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"85BBEAE208") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"16110193F34812E04E23FA1871F3E014") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"85BBEAE208";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"16110193F34812E04E23FA1871F3E014") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 191 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"85BBEAE208") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BD6AD594FB31559BFB6FF2175DFF4664") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"85BBEAE208";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BD6AD594FB31559BFB6FF2175DFF4664") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 192 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"85BBEAE208") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A40ECB65FA448E4B5FF5AE6D23182D24") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"85BBEAE208";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A40ECB65FA448E4B5FF5AE6D23182D24") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 193 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"85BBEAE208") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"11DE31A4F490F68D6F90D7317F9B0A17") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"85BBEAE208";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"11DE31A4F490F68D6F90D7317F9B0A17") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 194 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"85BBEAE208") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DFA0461E28D463536931B9FD5CBC3955") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"85BBEAE208";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DFA0461E28D463536931B9FD5CBC3955") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 195 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"85BBEAE208") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"655B0C2B627731F50AC880A5095DE25E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"85BBEAE208";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"655B0C2B627731F50AC880A5095DE25E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 196 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"85BBEAE208") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C6E077609B06F28FDB2BA77E6969915B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"85BBEAE208";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C6E077609B06F28FDB2BA77E6969915B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 197 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"85BBEAE208") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9E51079377B9705AAAA196A61DA3E530") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"85BBEAE208";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9E51079377B9705AAAA196A61DA3E530") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 198 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"85BBEAE208") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A09CB200FD93993FBA0062B045A8A5BF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"85BBEAE208";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A09CB200FD93993FBA0062B045A8A5BF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 199 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"85BBEAE208B7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"27721308E0575CD9A3DEB36EBB60883A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"85BBEAE208B7";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"27721308E0575CD9A3DEB36EBB60883A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 200 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"85BBEAE208B7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F99C930DAD872FE09E9E5E174B4732A3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"85BBEAE208B7";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F99C930DAD872FE09E9E5E174B4732A3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 201 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"85BBEAE208B7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D8B45523C875634427298747CF1F537C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"85BBEAE208B7";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D8B45523C875634427298747CF1F537C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 202 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"85BBEAE208B7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7C23A4D970845E380A9BFE443EBE8FE3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"85BBEAE208B7";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7C23A4D970845E380A9BFE443EBE8FE3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 203 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"85BBEAE208B7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"74A555E695900EAA4B1CEE531DFAF2D0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"85BBEAE208B7";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"74A555E695900EAA4B1CEE531DFAF2D0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 204 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"85BBEAE208B7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6036196AD2B5FC863203153BF58CA87A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"85BBEAE208B7";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6036196AD2B5FC863203153BF58CA87A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 205 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"85BBEAE208B7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"544B0889AD6A9B82802B103EA6C94028") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"85BBEAE208B7";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"544B0889AD6A9B82802B103EA6C94028") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 206 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"85BBEAE208B7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"69CD7961B7AE3BE263EDC2C94A419DB8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"85BBEAE208B7";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"69CD7961B7AE3BE263EDC2C94A419DB8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 207 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"85BBEAE208B7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"443F98E74DCC0A726669252BABB03876") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"85BBEAE208B7";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"443F98E74DCC0A726669252BABB03876") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 208 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"85BBEAE208B7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"754C5D7DB253FEEAC2DDE2BEAD15DB36") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"85BBEAE208B7";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"754C5D7DB253FEEAC2DDE2BEAD15DB36") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 209 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"85BBEAE208B7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"86D03C8AA0DF7AB462998DEE8E93E439") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"85BBEAE208B7";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"86D03C8AA0DF7AB462998DEE8E93E439") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 210 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"85BBEAE208B7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BDCCD7438F280DF28E312390B6B3B68D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"85BBEAE208B7";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BDCCD7438F280DF28E312390B6B3B68D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 211 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"85BBEAE208B7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"461D98DB8065108555B56576139E6361") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"85BBEAE208B7";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"461D98DB8065108555B56576139E6361") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 212 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"85BBEAE208B7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CC7171626A9F00FF933F69ED832436FE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"85BBEAE208B7";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CC7171626A9F00FF933F69ED832436FE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 213 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"85BBEAE208B7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FDAB246A6A2E4F587BAF7630528F9278") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"85BBEAE208B7";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FDAB246A6A2E4F587BAF7630528F9278") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 214 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"85BBEAE208B7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7877FB62F655964E771BADBB28CA3574") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"85BBEAE208B7";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7877FB62F655964E771BADBB28CA3574") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 215 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"85BBEAE208B7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C8F6A03F5D56D0C94F3DECDD21617DAA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"85BBEAE208B7";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C8F6A03F5D56D0C94F3DECDD21617DAA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 216 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"85BBEAE208B7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"76F098EA6E8612C9B7408B4F1826F640") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"85BBEAE208B7";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"76F098EA6E8612C9B7408B4F1826F640") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 217 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"85BBEAE208B7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"495E6C80A5864CE211E738A64584D8FD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"85BBEAE208B7";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"495E6C80A5864CE211E738A64584D8FD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 218 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"85BBEAE208B7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D12914AA859617106DF92E789E0AAB2D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"85BBEAE208B7";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D12914AA859617106DF92E789E0AAB2D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 219 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"85BBEAE208B7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AD1FF59F6128DCBF708B39EF80797E9A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"85BBEAE208B7";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AD1FF59F6128DCBF708B39EF80797E9A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 220 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"85BBEAE208B7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"ADFFA544798CE9BB41907B0C0802B8C8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"85BBEAE208B7";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"ADFFA544798CE9BB41907B0C0802B8C8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 221 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"85BBEAE208B7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7E063492CD8AB2C96BD2C31CEA8E7047") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"85BBEAE208B7";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7E063492CD8AB2C96BD2C31CEA8E7047") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 222 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"85BBEAE208B7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B8133488CDC552AAC34D757EEB1247C5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"85BBEAE208B7";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B8133488CDC552AAC34D757EEB1247C5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 223 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"85BBEAE208B7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3E0A6C6470B364B120975ADACC097953") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"85BBEAE208B7";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3E0A6C6470B364B120975ADACC097953") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 224 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"85BBEAE208B7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9571B86378CA23CA95DB52D5E005DF23") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"85BBEAE208B7";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9571B86378CA23CA95DB52D5E005DF23") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 225 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"85BBEAE208B7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8C15A69279BFF81A31410EAF9EE2B463") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"85BBEAE208B7";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8C15A69279BFF81A31410EAF9EE2B463") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 226 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"85BBEAE208B7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"39C55C53776B80DC012477F3C2619350") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"85BBEAE208B7";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"39C55C53776B80DC012477F3C2619350") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 227 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"85BBEAE208B7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F7BB2BE9AB2F15020785193FE146A012") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"85BBEAE208B7";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F7BB2BE9AB2F15020785193FE146A012") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 228 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"85BBEAE208B7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4D4061DCE18C47A4647C2067B4A77B19") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"85BBEAE208B7";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4D4061DCE18C47A4647C2067B4A77B19") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 229 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"85BBEAE208B7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EEFB1A9718FD84DEB59F07BCD493081C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"85BBEAE208B7";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EEFB1A9718FD84DEB59F07BCD493081C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 230 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"85BBEAE208B7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B64A6A64F442060BC4153664A0597C77") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"85BBEAE208B7";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B64A6A64F442060BC4153664A0597C77") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 231 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"85BBEAE208B7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8887DFF77E68EF6ED4B4C272F8523CF8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"85BBEAE208B7";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8887DFF77E68EF6ED4B4C272F8523CF8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 232 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"85BBEAE208B70D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2D307A9627796451E9DCAE28F8B3D0E6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"85BBEAE208B70D";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2D307A9627796451E9DCAE28F8B3D0E6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 233 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"85BBEAE208B70D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F3DEFA936AA91768D49C435108946A7F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"85BBEAE208B70D";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F3DEFA936AA91768D49C435108946A7F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 234 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"85BBEAE208B70D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D2F63CBD0F5B5BCC6D2B9A018CCC0BA0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"85BBEAE208B70D";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D2F63CBD0F5B5BCC6D2B9A018CCC0BA0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 235 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"85BBEAE208B70D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7661CD47B7AA66B04099E3027D6DD73F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"85BBEAE208B70D";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7661CD47B7AA66B04099E3027D6DD73F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 236 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"85BBEAE208B70D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7EE73C7852BE3622011EF3155E29AA0C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"85BBEAE208B70D";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7EE73C7852BE3622011EF3155E29AA0C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 237 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"85BBEAE208B70D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6A7470F4159BC40E7801087DB65FF0A6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"85BBEAE208B70D";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6A7470F4159BC40E7801087DB65FF0A6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 238 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"85BBEAE208B70D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5E0961176A44A30ACA290D78E51A18F4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"85BBEAE208B70D";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5E0961176A44A30ACA290D78E51A18F4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 239 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"85BBEAE208B70D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"638F10FF7080036A29EFDF8F0992C564") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"85BBEAE208B70D";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"638F10FF7080036A29EFDF8F0992C564") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 240 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"85BBEAE208B70D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4E7DF1798AE232FA2C6B386DE86360AA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"85BBEAE208B70D";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4E7DF1798AE232FA2C6B386DE86360AA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 241 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"85BBEAE208B70D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7F0E34E3757DC66288DFFFF8EEC683EA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"85BBEAE208B70D";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7F0E34E3757DC66288DFFFF8EEC683EA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 242 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"85BBEAE208B70D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8C92551467F1423C289B90A8CD40BCE5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"85BBEAE208B70D";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8C92551467F1423C289B90A8CD40BCE5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 243 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"85BBEAE208B70D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B78EBEDD4806357AC4333ED6F560EE51") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"85BBEAE208B70D";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B78EBEDD4806357AC4333ED6F560EE51") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 244 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"85BBEAE208B70D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4C5FF145474B280D1FB77830504D3BBD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"85BBEAE208B70D";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4C5FF145474B280D1FB77830504D3BBD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 245 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"85BBEAE208B70D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C63318FCADB13877D93D74ABC0F76E22") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"85BBEAE208B70D";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C63318FCADB13877D93D74ABC0F76E22") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 246 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"85BBEAE208B70D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F7E94DF4AD0077D031AD6B76115CCAA4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"85BBEAE208B70D";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F7E94DF4AD0077D031AD6B76115CCAA4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 247 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"85BBEAE208B70D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"723592FC317BAEC63D19B0FD6B196DA8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"85BBEAE208B70D";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"723592FC317BAEC63D19B0FD6B196DA8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 248 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"85BBEAE208B70D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C2B4C9A19A78E841053FF19B62B22576") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"85BBEAE208B70D";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C2B4C9A19A78E841053FF19B62B22576") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 249 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"85BBEAE208B70D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7CB2F174A9A82A41FD4296095BF5AE9C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"85BBEAE208B70D";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7CB2F174A9A82A41FD4296095BF5AE9C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 250 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"85BBEAE208B70D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"431C051E62A8746A5BE525E006578021") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"85BBEAE208B70D";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"431C051E62A8746A5BE525E006578021") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 251 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"85BBEAE208B70D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DB6B7D3442B82F9827FB333EDDD9F3F1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"85BBEAE208B70D";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DB6B7D3442B82F9827FB333EDDD9F3F1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 252 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"85BBEAE208B70D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A75D9C01A606E4373A8924A9C3AA2646") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"85BBEAE208B70D";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A75D9C01A606E4373A8924A9C3AA2646") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 253 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"85BBEAE208B70D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A7BDCCDABEA2D1330B92664A4BD1E014") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"85BBEAE208B70D";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A7BDCCDABEA2D1330B92664A4BD1E014") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 254 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"85BBEAE208B70D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"74445D0C0AA48A4121D0DE5AA95D289B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"85BBEAE208B70D";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"74445D0C0AA48A4121D0DE5AA95D289B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 255 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"85BBEAE208B70D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B2515D160AEB6A22894F6838A8C11F19") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"85BBEAE208B70D";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B2515D160AEB6A22894F6838A8C11F19") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 256 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"85BBEAE208B70D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"344805FAB79D5C396A95479C8FDA218F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"85BBEAE208B70D";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"344805FAB79D5C396A95479C8FDA218F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 257 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"85BBEAE208B70D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9F33D1FDBFE41B42DFD94F93A3D687FF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"85BBEAE208B70D";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9F33D1FDBFE41B42DFD94F93A3D687FF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 258 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"85BBEAE208B70D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8657CF0CBE91C0927B4313E9DD31ECBF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"85BBEAE208B70D";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8657CF0CBE91C0927B4313E9DD31ECBF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 259 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"85BBEAE208B70D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"338735CDB045B8544B266AB581B2CB8C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"85BBEAE208B70D";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"338735CDB045B8544B266AB581B2CB8C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 260 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"85BBEAE208B70D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FDF942776C012D8A4D870479A295F8CE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"85BBEAE208B70D";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FDF942776C012D8A4D870479A295F8CE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 261 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"85BBEAE208B70D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4702084226A27F2C2E7E3D21F77423C5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"85BBEAE208B70D";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4702084226A27F2C2E7E3D21F77423C5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 262 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"85BBEAE208B70D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E4B97309DFD3BC56FF9D1AFA974050C0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"85BBEAE208B70D";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E4B97309DFD3BC56FF9D1AFA974050C0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 263 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"85BBEAE208B70D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BC0803FA336C3E838E172B22E38A24AB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"85BBEAE208B70D";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BC0803FA336C3E838E172B22E38A24AB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 264 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"85BBEAE208B70D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"82C5B669B946D7E69EB6DF34BB816424") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"85BBEAE208B70D";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"82C5B669B946D7E69EB6DF34BB816424") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 265 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"85BBEAE208B70D61") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D31D1AEA2FBAD8B817EFE1DBC8168988") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"85BBEAE208B70D61";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D31D1AEA2FBAD8B817EFE1DBC8168988") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 266 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"85BBEAE208B70D61") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0DF39AEF626AAB812AAF0CA238313311") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"85BBEAE208B70D61";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0DF39AEF626AAB812AAF0CA238313311") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 267 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"85BBEAE208B70D61") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2CDB5CC10798E7259318D5F2BC6952CE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"85BBEAE208B70D61";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2CDB5CC10798E7259318D5F2BC6952CE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 268 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"85BBEAE208B70D61") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"884CAD3BBF69DA59BEAAACF14DC88E51") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"85BBEAE208B70D61";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"884CAD3BBF69DA59BEAAACF14DC88E51") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 269 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"85BBEAE208B70D61") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"80CA5C045A7D8ACBFF2DBCE66E8CF362") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"85BBEAE208B70D61";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"80CA5C045A7D8ACBFF2DBCE66E8CF362") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 270 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"85BBEAE208B70D61") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"945910881D5878E78632478E86FAA9C8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"85BBEAE208B70D61";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"945910881D5878E78632478E86FAA9C8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 271 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"85BBEAE208B70D61") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A024016B62871FE3341A428BD5BF419A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"85BBEAE208B70D61";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A024016B62871FE3341A428BD5BF419A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 272 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"85BBEAE208B70D61") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9DA270837843BF83D7DC907C39379C0A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"85BBEAE208B70D61";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9DA270837843BF83D7DC907C39379C0A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 273 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"85BBEAE208B70D61") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B050910582218E13D258779ED8C639C4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"85BBEAE208B70D61";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B050910582218E13D258779ED8C639C4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 274 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"85BBEAE208B70D61") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8123549F7DBE7A8B76ECB00BDE63DA84") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"85BBEAE208B70D61";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8123549F7DBE7A8B76ECB00BDE63DA84") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 275 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"85BBEAE208B70D61") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"72BF35686F32FED5D6A8DF5BFDE5E58B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"85BBEAE208B70D61";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"72BF35686F32FED5D6A8DF5BFDE5E58B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 276 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"85BBEAE208B70D61") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"49A3DEA140C589933A007125C5C5B73F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"85BBEAE208B70D61";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"49A3DEA140C589933A007125C5C5B73F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 277 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"85BBEAE208B70D61") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B27291394F8894E4E18437C360E862D3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"85BBEAE208B70D61";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B27291394F8894E4E18437C360E862D3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 278 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"85BBEAE208B70D61") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"381E7880A572849E270E3B58F052374C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"85BBEAE208B70D61";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"381E7880A572849E270E3B58F052374C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 279 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"85BBEAE208B70D61") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"09C42D88A5C3CB39CF9E248521F993CA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"85BBEAE208B70D61";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"09C42D88A5C3CB39CF9E248521F993CA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 280 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"85BBEAE208B70D61") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8C18F28039B8122FC32AFF0E5BBC34C6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"85BBEAE208B70D61";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8C18F28039B8122FC32AFF0E5BBC34C6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 281 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"85BBEAE208B70D61") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3C99A9DD92BB54A8FB0CBE6852177C18") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"85BBEAE208B70D61";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3C99A9DD92BB54A8FB0CBE6852177C18") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 282 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"85BBEAE208B70D61") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"829F9108A16B96A80371D9FA6B50F7F2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"85BBEAE208B70D61";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"829F9108A16B96A80371D9FA6B50F7F2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 283 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"85BBEAE208B70D61") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BD3165626A6BC883A5D66A1336F2D94F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"85BBEAE208B70D61";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BD3165626A6BC883A5D66A1336F2D94F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 284 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"85BBEAE208B70D61") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"25461D484A7B9371D9C87CCDED7CAA9F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"85BBEAE208B70D61";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"25461D484A7B9371D9C87CCDED7CAA9F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 285 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"85BBEAE208B70D61") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5970FC7DAEC558DEC4BA6B5AF30F7F28") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"85BBEAE208B70D61";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5970FC7DAEC558DEC4BA6B5AF30F7F28") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 286 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"85BBEAE208B70D61") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5990ACA6B6616DDAF5A129B97B74B97A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"85BBEAE208B70D61";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5990ACA6B6616DDAF5A129B97B74B97A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 287 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"85BBEAE208B70D61") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8A693D70026736A8DFE391A999F871F5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"85BBEAE208B70D61";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8A693D70026736A8DFE391A999F871F5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 288 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"85BBEAE208B70D61") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4C7C3D6A0228D6CB777C27CB98644677") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"85BBEAE208B70D61";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4C7C3D6A0228D6CB777C27CB98644677") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 289 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"85BBEAE208B70D61") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CA656586BF5EE0D094A6086FBF7F78E1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"85BBEAE208B70D61";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CA656586BF5EE0D094A6086FBF7F78E1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 290 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"85BBEAE208B70D61") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"611EB181B727A7AB21EA00609373DE91") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"85BBEAE208B70D61";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"611EB181B727A7AB21EA00609373DE91") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 291 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"85BBEAE208B70D61") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"787AAF70B6527C7B85705C1AED94B5D1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"85BBEAE208B70D61";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"787AAF70B6527C7B85705C1AED94B5D1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 292 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"85BBEAE208B70D61") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CDAA55B1B88604BDB5152546B11792E2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"85BBEAE208B70D61";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CDAA55B1B88604BDB5152546B11792E2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 293 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"85BBEAE208B70D61") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"03D4220B64C29163B3B44B8A9230A1A0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"85BBEAE208B70D61";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"03D4220B64C29163B3B44B8A9230A1A0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 294 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"85BBEAE208B70D61") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B92F683E2E61C3C5D04D72D2C7D17AAB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"85BBEAE208B70D61";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B92F683E2E61C3C5D04D72D2C7D17AAB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 295 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"85BBEAE208B70D61") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1A941375D71000BF01AE5509A7E509AE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"85BBEAE208B70D61";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1A941375D71000BF01AE5509A7E509AE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 296 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"85BBEAE208B70D61") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"422563863BAF826A702464D1D32F7DC5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"85BBEAE208B70D61";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"422563863BAF826A702464D1D32F7DC5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 297 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"85BBEAE208B70D61") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7CE8D615B1856B0F608590C78B243D4A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"85BBEAE208B70D61";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7CE8D615B1856B0F608590C78B243D4A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 298 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"85BBEAE208B70D615C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1DD08BB76F55C61540509898E91351F7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"85BBEAE208B70D615C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1DD08BB76F55C61540509898E91351F7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 299 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"85BBEAE208B70D615C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C33E0BB22285B52C7D1075E11934EB6E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"85BBEAE208B70D615C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C33E0BB22285B52C7D1075E11934EB6E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 300 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"85BBEAE208B70D615C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E216CD9C4777F988C4A7ACB19D6C8AB1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"85BBEAE208B70D615C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E216CD9C4777F988C4A7ACB19D6C8AB1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 301 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"85BBEAE208B70D615C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"46813C66FF86C4F4E915D5B26CCD562E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"85BBEAE208B70D615C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"46813C66FF86C4F4E915D5B26CCD562E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 302 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"85BBEAE208B70D615C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4E07CD591A929466A892C5A54F892B1D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"85BBEAE208B70D615C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4E07CD591A929466A892C5A54F892B1D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 303 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"85BBEAE208B70D615C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5A9481D55DB7664AD18D3ECDA7FF71B7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"85BBEAE208B70D615C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5A9481D55DB7664AD18D3ECDA7FF71B7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 304 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"85BBEAE208B70D615C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6EE990362268014E63A53BC8F4BA99E5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"85BBEAE208B70D615C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6EE990362268014E63A53BC8F4BA99E5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 305 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"85BBEAE208B70D615C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"536FE1DE38ACA12E8063E93F18324475") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"85BBEAE208B70D615C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"536FE1DE38ACA12E8063E93F18324475") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 306 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"85BBEAE208B70D615C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7E9D0058C2CE90BE85E70EDDF9C3E1BB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"85BBEAE208B70D615C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7E9D0058C2CE90BE85E70EDDF9C3E1BB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 307 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"85BBEAE208B70D615C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4FEEC5C23D5164262153C948FF6602FB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"85BBEAE208B70D615C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4FEEC5C23D5164262153C948FF6602FB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 308 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"85BBEAE208B70D615C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BC72A4352FDDE0788117A618DCE03DF4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"85BBEAE208B70D615C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BC72A4352FDDE0788117A618DCE03DF4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 309 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"85BBEAE208B70D615C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"876E4FFC002A973E6DBF0866E4C06F40") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"85BBEAE208B70D615C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"876E4FFC002A973E6DBF0866E4C06F40") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 310 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"85BBEAE208B70D615C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7CBF00640F678A49B63B4E8041EDBAAC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"85BBEAE208B70D615C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7CBF00640F678A49B63B4E8041EDBAAC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 311 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"85BBEAE208B70D615C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F6D3E9DDE59D9A3370B1421BD157EF33") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"85BBEAE208B70D615C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F6D3E9DDE59D9A3370B1421BD157EF33") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 312 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"85BBEAE208B70D615C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C709BCD5E52CD59498215DC600FC4BB5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"85BBEAE208B70D615C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C709BCD5E52CD59498215DC600FC4BB5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 313 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"85BBEAE208B70D615C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"42D563DD79570C829495864D7AB9ECB9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"85BBEAE208B70D615C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"42D563DD79570C829495864D7AB9ECB9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 314 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"85BBEAE208B70D615C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F2543880D2544A05ACB3C72B7312A467") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"85BBEAE208B70D615C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F2543880D2544A05ACB3C72B7312A467") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 315 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"85BBEAE208B70D615C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4C520055E184880554CEA0B94A552F8D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"85BBEAE208B70D615C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4C520055E184880554CEA0B94A552F8D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 316 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"85BBEAE208B70D615C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"73FCF43F2A84D62EF269135017F70130") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"85BBEAE208B70D615C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"73FCF43F2A84D62EF269135017F70130") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 317 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"85BBEAE208B70D615C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EB8B8C150A948DDC8E77058ECC7972E0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"85BBEAE208B70D615C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EB8B8C150A948DDC8E77058ECC7972E0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 318 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"85BBEAE208B70D615C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"97BD6D20EE2A467393051219D20AA757") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"85BBEAE208B70D615C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"97BD6D20EE2A467393051219D20AA757") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 319 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"85BBEAE208B70D615C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"975D3DFBF68E7377A21E50FA5A716105") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"85BBEAE208B70D615C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"975D3DFBF68E7377A21E50FA5A716105") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 320 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"85BBEAE208B70D615C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"44A4AC2D42882805885CE8EAB8FDA98A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"85BBEAE208B70D615C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"44A4AC2D42882805885CE8EAB8FDA98A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 321 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"85BBEAE208B70D615C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"82B1AC3742C7C86620C35E88B9619E08") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"85BBEAE208B70D615C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"82B1AC3742C7C86620C35E88B9619E08") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 322 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"85BBEAE208B70D615C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"04A8F4DBFFB1FE7DC319712C9E7AA09E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"85BBEAE208B70D615C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"04A8F4DBFFB1FE7DC319712C9E7AA09E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 323 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"85BBEAE208B70D615C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AFD320DCF7C8B90676557923B27606EE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"85BBEAE208B70D615C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AFD320DCF7C8B90676557923B27606EE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 324 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"85BBEAE208B70D615C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B6B73E2DF6BD62D6D2CF2559CC916DAE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"85BBEAE208B70D615C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B6B73E2DF6BD62D6D2CF2559CC916DAE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 325 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"85BBEAE208B70D615C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0367C4ECF8691A10E2AA5C0590124A9D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"85BBEAE208B70D615C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0367C4ECF8691A10E2AA5C0590124A9D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 326 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"85BBEAE208B70D615C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CD19B356242D8FCEE40B32C9B33579DF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"85BBEAE208B70D615C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CD19B356242D8FCEE40B32C9B33579DF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 327 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"85BBEAE208B70D615C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"77E2F9636E8EDD6887F20B91E6D4A2D4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"85BBEAE208B70D615C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"77E2F9636E8EDD6887F20B91E6D4A2D4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 328 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"85BBEAE208B70D615C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D459822897FF1E1256112C4A86E0D1D1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"85BBEAE208B70D615C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D459822897FF1E1256112C4A86E0D1D1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 329 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"85BBEAE208B70D615C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8CE8F2DB7B409CC7279B1D92F22AA5BA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"85BBEAE208B70D615C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8CE8F2DB7B409CC7279B1D92F22AA5BA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 330 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"85BBEAE208B70D615C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B2254748F16A75A2373AE984AA21E535") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"85BBEAE208B70D615C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B2254748F16A75A2373AE984AA21E535") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 331 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"85BBEAE208B70D615C45") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"18BB0AA0E788B6E9C9E995BEDCA49A08") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"85BBEAE208B70D615C45";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"18BB0AA0E788B6E9C9E995BEDCA49A08") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 332 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"85BBEAE208B70D615C45") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C6558AA5AA58C5D0F4A978C72C832091") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"85BBEAE208B70D615C45";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C6558AA5AA58C5D0F4A978C72C832091") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 333 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"85BBEAE208B70D615C45") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E77D4C8BCFAA89744D1EA197A8DB414E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"85BBEAE208B70D615C45";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E77D4C8BCFAA89744D1EA197A8DB414E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 334 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"85BBEAE208B70D615C45") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"43EABD71775BB40860ACD894597A9DD1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"85BBEAE208B70D615C45";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"43EABD71775BB40860ACD894597A9DD1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 335 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"85BBEAE208B70D615C45") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4B6C4C4E924FE49A212BC8837A3EE0E2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"85BBEAE208B70D615C45";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4B6C4C4E924FE49A212BC8837A3EE0E2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 336 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"85BBEAE208B70D615C45") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5FFF00C2D56A16B6583433EB9248BA48") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"85BBEAE208B70D615C45";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5FFF00C2D56A16B6583433EB9248BA48") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 337 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"85BBEAE208B70D615C45") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6B821121AAB571B2EA1C36EEC10D521A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"85BBEAE208B70D615C45";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6B821121AAB571B2EA1C36EEC10D521A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 338 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"85BBEAE208B70D615C45") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"560460C9B071D1D209DAE4192D858F8A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"85BBEAE208B70D615C45";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"560460C9B071D1D209DAE4192D858F8A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 339 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"85BBEAE208B70D615C45") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7BF6814F4A13E0420C5E03FBCC742A44") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"85BBEAE208B70D615C45";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7BF6814F4A13E0420C5E03FBCC742A44") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 340 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"85BBEAE208B70D615C45") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4A8544D5B58C14DAA8EAC46ECAD1C904") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"85BBEAE208B70D615C45";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4A8544D5B58C14DAA8EAC46ECAD1C904") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 341 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"85BBEAE208B70D615C45") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B9192522A700908408AEAB3EE957F60B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"85BBEAE208B70D615C45";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B9192522A700908408AEAB3EE957F60B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 342 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"85BBEAE208B70D615C45") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8205CEEB88F7E7C2E4060540D177A4BF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"85BBEAE208B70D615C45";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8205CEEB88F7E7C2E4060540D177A4BF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 343 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"85BBEAE208B70D615C45") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"79D4817387BAFAB53F8243A6745A7153") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"85BBEAE208B70D615C45";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"79D4817387BAFAB53F8243A6745A7153") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 344 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"85BBEAE208B70D615C45") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F3B868CA6D40EACFF9084F3DE4E024CC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"85BBEAE208B70D615C45";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F3B868CA6D40EACFF9084F3DE4E024CC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 345 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"85BBEAE208B70D615C45") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C2623DC26DF1A568119850E0354B804A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"85BBEAE208B70D615C45";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C2623DC26DF1A568119850E0354B804A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 346 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"85BBEAE208B70D615C45") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"47BEE2CAF18A7C7E1D2C8B6B4F0E2746") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"85BBEAE208B70D615C45";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"47BEE2CAF18A7C7E1D2C8B6B4F0E2746") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 347 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"85BBEAE208B70D615C45") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F73FB9975A893AF9250ACA0D46A56F98") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"85BBEAE208B70D615C45";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F73FB9975A893AF9250ACA0D46A56F98") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 348 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"85BBEAE208B70D615C45") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"493981426959F8F9DD77AD9F7FE2E472") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"85BBEAE208B70D615C45";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"493981426959F8F9DD77AD9F7FE2E472") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 349 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"85BBEAE208B70D615C45") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"76977528A259A6D27BD01E762240CACF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"85BBEAE208B70D615C45";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"76977528A259A6D27BD01E762240CACF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 350 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"85BBEAE208B70D615C45") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EEE00D028249FD2007CE08A8F9CEB91F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"85BBEAE208B70D615C45";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EEE00D028249FD2007CE08A8F9CEB91F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 351 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"85BBEAE208B70D615C45") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"92D6EC3766F7368F1ABC1F3FE7BD6CA8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"85BBEAE208B70D615C45";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"92D6EC3766F7368F1ABC1F3FE7BD6CA8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 352 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"85BBEAE208B70D615C45") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9236BCEC7E53038B2BA75DDC6FC6AAFA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"85BBEAE208B70D615C45";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9236BCEC7E53038B2BA75DDC6FC6AAFA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 353 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"85BBEAE208B70D615C45") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"41CF2D3ACA5558F901E5E5CC8D4A6275") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"85BBEAE208B70D615C45";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"41CF2D3ACA5558F901E5E5CC8D4A6275") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 354 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"85BBEAE208B70D615C45") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"87DA2D20CA1AB89AA97A53AE8CD655F7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"85BBEAE208B70D615C45";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"87DA2D20CA1AB89AA97A53AE8CD655F7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 355 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"85BBEAE208B70D615C45") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"01C375CC776C8E814AA07C0AABCD6B61") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"85BBEAE208B70D615C45";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"01C375CC776C8E814AA07C0AABCD6B61") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 356 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"85BBEAE208B70D615C45") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AAB8A1CB7F15C9FAFFEC740587C1CD11") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"85BBEAE208B70D615C45";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AAB8A1CB7F15C9FAFFEC740587C1CD11") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 357 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"85BBEAE208B70D615C45") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B3DCBF3A7E60122A5B76287FF926A651") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"85BBEAE208B70D615C45";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B3DCBF3A7E60122A5B76287FF926A651") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 358 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"85BBEAE208B70D615C45") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"060C45FB70B46AEC6B135123A5A58162") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"85BBEAE208B70D615C45";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"060C45FB70B46AEC6B135123A5A58162") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 359 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"85BBEAE208B70D615C45") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C8723241ACF0FF326DB23FEF8682B220") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"85BBEAE208B70D615C45";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C8723241ACF0FF326DB23FEF8682B220") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 360 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"85BBEAE208B70D615C45") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"72897874E653AD940E4B06B7D363692B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"85BBEAE208B70D615C45";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"72897874E653AD940E4B06B7D363692B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 361 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"85BBEAE208B70D615C45") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D132033F1F226EEEDFA8216CB3571A2E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"85BBEAE208B70D615C45";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D132033F1F226EEEDFA8216CB3571A2E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 362 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"85BBEAE208B70D615C45") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"898373CCF39DEC3BAE2210B4C79D6E45") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"85BBEAE208B70D615C45";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"898373CCF39DEC3BAE2210B4C79D6E45") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 363 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"85BBEAE208B70D615C45") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B74EC65F79B7055EBE83E4A29F962ECA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"85BBEAE208B70D615C45";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B74EC65F79B7055EBE83E4A29F962ECA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 364 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"85BBEAE208B70D615C45F7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3D6EEA04D78181B3DC284AE97826A626") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"85BBEAE208B70D615C45F7";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3D6EEA04D78181B3DC284AE97826A626") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 365 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"85BBEAE208B70D615C45F7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E3806A019A51F28AE168A79088011CBF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"85BBEAE208B70D615C45F7";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E3806A019A51F28AE168A79088011CBF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 366 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"85BBEAE208B70D615C45F7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C2A8AC2FFFA3BE2E58DF7EC00C597D60") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"85BBEAE208B70D615C45F7";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C2A8AC2FFFA3BE2E58DF7EC00C597D60") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 367 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"85BBEAE208B70D615C45F7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"663F5DD547528352756D07C3FDF8A1FF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"85BBEAE208B70D615C45F7";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"663F5DD547528352756D07C3FDF8A1FF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 368 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"85BBEAE208B70D615C45F7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6EB9ACEAA246D3C034EA17D4DEBCDCCC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"85BBEAE208B70D615C45F7";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6EB9ACEAA246D3C034EA17D4DEBCDCCC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 369 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"85BBEAE208B70D615C45F7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7A2AE066E56321EC4DF5ECBC36CA8666") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"85BBEAE208B70D615C45F7";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7A2AE066E56321EC4DF5ECBC36CA8666") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 370 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"85BBEAE208B70D615C45F7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4E57F1859ABC46E8FFDDE9B9658F6E34") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"85BBEAE208B70D615C45F7";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4E57F1859ABC46E8FFDDE9B9658F6E34") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 371 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"85BBEAE208B70D615C45F7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"73D1806D8078E6881C1B3B4E8907B3A4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"85BBEAE208B70D615C45F7";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"73D1806D8078E6881C1B3B4E8907B3A4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 372 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"85BBEAE208B70D615C45F7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5E2361EB7A1AD718199FDCAC68F6166A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"85BBEAE208B70D615C45F7";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5E2361EB7A1AD718199FDCAC68F6166A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 373 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"85BBEAE208B70D615C45F7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6F50A47185852380BD2B1B396E53F52A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"85BBEAE208B70D615C45F7";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6F50A47185852380BD2B1B396E53F52A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 374 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"85BBEAE208B70D615C45F7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9CCCC5869709A7DE1D6F74694DD5CA25") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"85BBEAE208B70D615C45F7";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9CCCC5869709A7DE1D6F74694DD5CA25") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 375 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"85BBEAE208B70D615C45F7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A7D02E4FB8FED098F1C7DA1775F59891") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"85BBEAE208B70D615C45F7";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A7D02E4FB8FED098F1C7DA1775F59891") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 376 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"85BBEAE208B70D615C45F7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5C0161D7B7B3CDEF2A439CF1D0D84D7D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"85BBEAE208B70D615C45F7";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5C0161D7B7B3CDEF2A439CF1D0D84D7D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 377 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"85BBEAE208B70D615C45F7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D66D886E5D49DD95ECC9906A406218E2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"85BBEAE208B70D615C45F7";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D66D886E5D49DD95ECC9906A406218E2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 378 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"85BBEAE208B70D615C45F7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E7B7DD665DF8923204598FB791C9BC64") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"85BBEAE208B70D615C45F7";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E7B7DD665DF8923204598FB791C9BC64") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 379 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"85BBEAE208B70D615C45F7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"626B026EC1834B2408ED543CEB8C1B68") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"85BBEAE208B70D615C45F7";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"626B026EC1834B2408ED543CEB8C1B68") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 380 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"85BBEAE208B70D615C45F7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D2EA59336A800DA330CB155AE22753B6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"85BBEAE208B70D615C45F7";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D2EA59336A800DA330CB155AE22753B6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 381 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"85BBEAE208B70D615C45F7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6CEC61E65950CFA3C8B672C8DB60D85C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"85BBEAE208B70D615C45F7";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6CEC61E65950CFA3C8B672C8DB60D85C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 382 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"85BBEAE208B70D615C45F7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5342958C925091886E11C12186C2F6E1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"85BBEAE208B70D615C45F7";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5342958C925091886E11C12186C2F6E1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 383 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"85BBEAE208B70D615C45F7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CB35EDA6B240CA7A120FD7FF5D4C8531") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"85BBEAE208B70D615C45F7";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CB35EDA6B240CA7A120FD7FF5D4C8531") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 384 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"85BBEAE208B70D615C45F7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B7030C9356FE01D50F7DC068433F5086") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"85BBEAE208B70D615C45F7";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B7030C9356FE01D50F7DC068433F5086") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 385 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"85BBEAE208B70D615C45F7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B7E35C484E5A34D13E66828BCB4496D4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"85BBEAE208B70D615C45F7";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B7E35C484E5A34D13E66828BCB4496D4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 386 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"85BBEAE208B70D615C45F7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"641ACD9EFA5C6FA314243A9B29C85E5B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"85BBEAE208B70D615C45F7";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"641ACD9EFA5C6FA314243A9B29C85E5B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 387 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"85BBEAE208B70D615C45F7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A20FCD84FA138FC0BCBB8CF9285469D9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"85BBEAE208B70D615C45F7";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A20FCD84FA138FC0BCBB8CF9285469D9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 388 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"85BBEAE208B70D615C45F7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"241695684765B9DB5F61A35D0F4F574F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"85BBEAE208B70D615C45F7";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"241695684765B9DB5F61A35D0F4F574F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 389 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"85BBEAE208B70D615C45F7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8F6D416F4F1CFEA0EA2DAB522343F13F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"85BBEAE208B70D615C45F7";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8F6D416F4F1CFEA0EA2DAB522343F13F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 390 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"85BBEAE208B70D615C45F7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"96095F9E4E6925704EB7F7285DA49A7F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"85BBEAE208B70D615C45F7";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"96095F9E4E6925704EB7F7285DA49A7F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 391 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"85BBEAE208B70D615C45F7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"23D9A55F40BD5DB67ED28E740127BD4C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"85BBEAE208B70D615C45F7";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"23D9A55F40BD5DB67ED28E740127BD4C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 392 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"85BBEAE208B70D615C45F7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EDA7D2E59CF9C8687873E0B822008E0E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"85BBEAE208B70D615C45F7";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EDA7D2E59CF9C8687873E0B822008E0E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 393 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"85BBEAE208B70D615C45F7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"575C98D0D65A9ACE1B8AD9E077E15505") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"85BBEAE208B70D615C45F7";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"575C98D0D65A9ACE1B8AD9E077E15505") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 394 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"85BBEAE208B70D615C45F7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F4E7E39B2F2B59B4CA69FE3B17D52600") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"85BBEAE208B70D615C45F7";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F4E7E39B2F2B59B4CA69FE3B17D52600") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 395 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"85BBEAE208B70D615C45F7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AC569368C394DB61BBE3CFE3631F526B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"85BBEAE208B70D615C45F7";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AC569368C394DB61BBE3CFE3631F526B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 396 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"85BBEAE208B70D615C45F7") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"929B26FB49BE3204AB423BF53B1412E4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"85BBEAE208B70D615C45F7";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"929B26FB49BE3204AB423BF53B1412E4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 397 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"85BBEAE208B70D615C45F7BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4CE614EBAB68006E5DC33478A9F0DC88") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"85BBEAE208B70D615C45F7BC";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4CE614EBAB68006E5DC33478A9F0DC88") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 398 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"85BBEAE208B70D615C45F7BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"920894EEE6B873576083D90159D76611") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"85BBEAE208B70D615C45F7BC";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"920894EEE6B873576083D90159D76611") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 399 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"85BBEAE208B70D615C45F7BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B32052C0834A3FF3D9340051DD8F07CE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"85BBEAE208B70D615C45F7BC";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B32052C0834A3FF3D9340051DD8F07CE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 400 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"85BBEAE208B70D615C45F7BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"17B7A33A3BBB028FF48679522C2EDB51") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"85BBEAE208B70D615C45F7BC";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"17B7A33A3BBB028FF48679522C2EDB51") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 401 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"85BBEAE208B70D615C45F7BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1F315205DEAF521DB50169450F6AA662") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"85BBEAE208B70D615C45F7BC";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1F315205DEAF521DB50169450F6AA662") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 402 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"85BBEAE208B70D615C45F7BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0BA21E89998AA031CC1E922DE71CFCC8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"85BBEAE208B70D615C45F7BC";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0BA21E89998AA031CC1E922DE71CFCC8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 403 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"85BBEAE208B70D615C45F7BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3FDF0F6AE655C7357E369728B459149A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"85BBEAE208B70D615C45F7BC";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3FDF0F6AE655C7357E369728B459149A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 404 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"85BBEAE208B70D615C45F7BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"02597E82FC9167559DF045DF58D1C90A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"85BBEAE208B70D615C45F7BC";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"02597E82FC9167559DF045DF58D1C90A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 405 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"85BBEAE208B70D615C45F7BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2FAB9F0406F356C59874A23DB9206CC4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"85BBEAE208B70D615C45F7BC";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2FAB9F0406F356C59874A23DB9206CC4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 406 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"85BBEAE208B70D615C45F7BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1ED85A9EF96CA25D3CC065A8BF858F84") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"85BBEAE208B70D615C45F7BC";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1ED85A9EF96CA25D3CC065A8BF858F84") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 407 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"85BBEAE208B70D615C45F7BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"ED443B69EBE026039C840AF89C03B08B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"85BBEAE208B70D615C45F7BC";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"ED443B69EBE026039C840AF89C03B08B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 408 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"85BBEAE208B70D615C45F7BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D658D0A0C4175145702CA486A423E23F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"85BBEAE208B70D615C45F7BC";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D658D0A0C4175145702CA486A423E23F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 409 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"85BBEAE208B70D615C45F7BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2D899F38CB5A4C32ABA8E260010E37D3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"85BBEAE208B70D615C45F7BC";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2D899F38CB5A4C32ABA8E260010E37D3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 410 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"85BBEAE208B70D615C45F7BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A7E5768121A05C486D22EEFB91B4624C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"85BBEAE208B70D615C45F7BC";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A7E5768121A05C486D22EEFB91B4624C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 411 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"85BBEAE208B70D615C45F7BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"963F2389211113EF85B2F126401FC6CA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"85BBEAE208B70D615C45F7BC";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"963F2389211113EF85B2F126401FC6CA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 412 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"85BBEAE208B70D615C45F7BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"13E3FC81BD6ACAF989062AAD3A5A61C6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"85BBEAE208B70D615C45F7BC";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"13E3FC81BD6ACAF989062AAD3A5A61C6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 413 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"85BBEAE208B70D615C45F7BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A362A7DC16698C7EB1206BCB33F12918") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"85BBEAE208B70D615C45F7BC";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A362A7DC16698C7EB1206BCB33F12918") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 414 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"85BBEAE208B70D615C45F7BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1D649F0925B94E7E495D0C590AB6A2F2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"85BBEAE208B70D615C45F7BC";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1D649F0925B94E7E495D0C590AB6A2F2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 415 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"85BBEAE208B70D615C45F7BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"22CA6B63EEB91055EFFABFB057148C4F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"85BBEAE208B70D615C45F7BC";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"22CA6B63EEB91055EFFABFB057148C4F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 416 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"85BBEAE208B70D615C45F7BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BABD1349CEA94BA793E4A96E8C9AFF9F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"85BBEAE208B70D615C45F7BC";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BABD1349CEA94BA793E4A96E8C9AFF9F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 417 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"85BBEAE208B70D615C45F7BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C68BF27C2A1780088E96BEF992E92A28") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"85BBEAE208B70D615C45F7BC";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C68BF27C2A1780088E96BEF992E92A28") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 418 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"85BBEAE208B70D615C45F7BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C66BA2A732B3B50CBF8DFC1A1A92EC7A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"85BBEAE208B70D615C45F7BC";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C66BA2A732B3B50CBF8DFC1A1A92EC7A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 419 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"85BBEAE208B70D615C45F7BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1592337186B5EE7E95CF440AF81E24F5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"85BBEAE208B70D615C45F7BC";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1592337186B5EE7E95CF440AF81E24F5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 420 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"85BBEAE208B70D615C45F7BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D387336B86FA0E1D3D50F268F9821377") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"85BBEAE208B70D615C45F7BC";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D387336B86FA0E1D3D50F268F9821377") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 421 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"85BBEAE208B70D615C45F7BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"559E6B873B8C3806DE8ADDCCDE992DE1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"85BBEAE208B70D615C45F7BC";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"559E6B873B8C3806DE8ADDCCDE992DE1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 422 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"85BBEAE208B70D615C45F7BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FEE5BF8033F57F7D6BC6D5C3F2958B91") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"85BBEAE208B70D615C45F7BC";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FEE5BF8033F57F7D6BC6D5C3F2958B91") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 423 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"85BBEAE208B70D615C45F7BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E781A1713280A4ADCF5C89B98C72E0D1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"85BBEAE208B70D615C45F7BC";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E781A1713280A4ADCF5C89B98C72E0D1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 424 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"85BBEAE208B70D615C45F7BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"52515BB03C54DC6BFF39F0E5D0F1C7E2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"85BBEAE208B70D615C45F7BC";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"52515BB03C54DC6BFF39F0E5D0F1C7E2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 425 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"85BBEAE208B70D615C45F7BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9C2F2C0AE01049B5F9989E29F3D6F4A0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"85BBEAE208B70D615C45F7BC";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9C2F2C0AE01049B5F9989E29F3D6F4A0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 426 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"85BBEAE208B70D615C45F7BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"26D4663FAAB31B139A61A771A6372FAB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"85BBEAE208B70D615C45F7BC";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"26D4663FAAB31B139A61A771A6372FAB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 427 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"85BBEAE208B70D615C45F7BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"856F1D7453C2D8694B8280AAC6035CAE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"85BBEAE208B70D615C45F7BC";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"856F1D7453C2D8694B8280AAC6035CAE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 428 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"85BBEAE208B70D615C45F7BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DDDE6D87BF7D5ABC3A08B172B2C928C5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"85BBEAE208B70D615C45F7BC";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DDDE6D87BF7D5ABC3A08B172B2C928C5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 429 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"85BBEAE208B70D615C45F7BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E313D8143557B3D92AA94564EAC2684A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"85BBEAE208B70D615C45F7BC";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E313D8143557B3D92AA94564EAC2684A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 430 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"85BBEAE208B70D615C45F7BC62") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E037C054CB485C4E9166BA07497BFB8E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"85BBEAE208B70D615C45F7BC62";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E037C054CB485C4E9166BA07497BFB8E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 431 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"85BBEAE208B70D615C45F7BC62") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3ED9405186982F77AC26577EB95C4117") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"85BBEAE208B70D615C45F7BC62";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3ED9405186982F77AC26577EB95C4117") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 432 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"85BBEAE208B70D615C45F7BC62") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1FF1867FE36A63D315918E2E3D0420C8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"85BBEAE208B70D615C45F7BC62";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1FF1867FE36A63D315918E2E3D0420C8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 433 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"85BBEAE208B70D615C45F7BC62") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BB6677855B9B5EAF3823F72DCCA5FC57") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"85BBEAE208B70D615C45F7BC62";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BB6677855B9B5EAF3823F72DCCA5FC57") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 434 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"85BBEAE208B70D615C45F7BC62") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B3E086BABE8F0E3D79A4E73AEFE18164") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"85BBEAE208B70D615C45F7BC62";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B3E086BABE8F0E3D79A4E73AEFE18164") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 435 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"85BBEAE208B70D615C45F7BC62") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A773CA36F9AAFC1100BB1C520797DBCE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"85BBEAE208B70D615C45F7BC62";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A773CA36F9AAFC1100BB1C520797DBCE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 436 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"85BBEAE208B70D615C45F7BC62") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"930EDBD586759B15B293195754D2339C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"85BBEAE208B70D615C45F7BC62";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"930EDBD586759B15B293195754D2339C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 437 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"85BBEAE208B70D615C45F7BC62") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AE88AA3D9CB13B755155CBA0B85AEE0C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"85BBEAE208B70D615C45F7BC62";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AE88AA3D9CB13B755155CBA0B85AEE0C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 438 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"85BBEAE208B70D615C45F7BC62") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"837A4BBB66D30AE554D12C4259AB4BC2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"85BBEAE208B70D615C45F7BC62";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"837A4BBB66D30AE554D12C4259AB4BC2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 439 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"85BBEAE208B70D615C45F7BC62") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B2098E21994CFE7DF065EBD75F0EA882") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"85BBEAE208B70D615C45F7BC62";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B2098E21994CFE7DF065EBD75F0EA882") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 440 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"85BBEAE208B70D615C45F7BC62") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4195EFD68BC07A23502184877C88978D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"85BBEAE208B70D615C45F7BC62";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4195EFD68BC07A23502184877C88978D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 441 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"85BBEAE208B70D615C45F7BC62") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7A89041FA4370D65BC892AF944A8C539") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"85BBEAE208B70D615C45F7BC62";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7A89041FA4370D65BC892AF944A8C539") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 442 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"85BBEAE208B70D615C45F7BC62") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"81584B87AB7A1012670D6C1FE18510D5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"85BBEAE208B70D615C45F7BC62";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"81584B87AB7A1012670D6C1FE18510D5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 443 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"85BBEAE208B70D615C45F7BC62") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0B34A23E41800068A1876084713F454A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"85BBEAE208B70D615C45F7BC62";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0B34A23E41800068A1876084713F454A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 444 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"85BBEAE208B70D615C45F7BC62") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3AEEF73641314FCF49177F59A094E1CC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"85BBEAE208B70D615C45F7BC62";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3AEEF73641314FCF49177F59A094E1CC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 445 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"85BBEAE208B70D615C45F7BC62") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BF32283EDD4A96D945A3A4D2DAD146C0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"85BBEAE208B70D615C45F7BC62";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BF32283EDD4A96D945A3A4D2DAD146C0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 446 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"85BBEAE208B70D615C45F7BC62") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0FB373637649D05E7D85E5B4D37A0E1E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"85BBEAE208B70D615C45F7BC62";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0FB373637649D05E7D85E5B4D37A0E1E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 447 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"85BBEAE208B70D615C45F7BC62") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B1B54BB64599125E85F88226EA3D85F4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"85BBEAE208B70D615C45F7BC62";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B1B54BB64599125E85F88226EA3D85F4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 448 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"85BBEAE208B70D615C45F7BC62") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8E1BBFDC8E994C75235F31CFB79FAB49") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"85BBEAE208B70D615C45F7BC62";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8E1BBFDC8E994C75235F31CFB79FAB49") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 449 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"85BBEAE208B70D615C45F7BC62") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"166CC7F6AE8917875F4127116C11D899") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"85BBEAE208B70D615C45F7BC62";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"166CC7F6AE8917875F4127116C11D899") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 450 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"85BBEAE208B70D615C45F7BC62") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6A5A26C34A37DC284233308672620D2E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"85BBEAE208B70D615C45F7BC62";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6A5A26C34A37DC284233308672620D2E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 451 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"85BBEAE208B70D615C45F7BC62") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6ABA76185293E92C73287265FA19CB7C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"85BBEAE208B70D615C45F7BC62";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6ABA76185293E92C73287265FA19CB7C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 452 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"85BBEAE208B70D615C45F7BC62") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B943E7CEE695B25E596ACA75189503F3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"85BBEAE208B70D615C45F7BC62";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B943E7CEE695B25E596ACA75189503F3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 453 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"85BBEAE208B70D615C45F7BC62") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7F56E7D4E6DA523DF1F57C1719093471") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"85BBEAE208B70D615C45F7BC62";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7F56E7D4E6DA523DF1F57C1719093471") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 454 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"85BBEAE208B70D615C45F7BC62") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F94FBF385BAC6426122F53B33E120AE7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"85BBEAE208B70D615C45F7BC62";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F94FBF385BAC6426122F53B33E120AE7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 455 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"85BBEAE208B70D615C45F7BC62") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"52346B3F53D5235DA7635BBC121EAC97") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"85BBEAE208B70D615C45F7BC62";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"52346B3F53D5235DA7635BBC121EAC97") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 456 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"85BBEAE208B70D615C45F7BC62") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4B5075CE52A0F88D03F907C66CF9C7D7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"85BBEAE208B70D615C45F7BC62";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4B5075CE52A0F88D03F907C66CF9C7D7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 457 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"85BBEAE208B70D615C45F7BC62") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FE808F0F5C74804B339C7E9A307AE0E4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"85BBEAE208B70D615C45F7BC62";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FE808F0F5C74804B339C7E9A307AE0E4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 458 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"85BBEAE208B70D615C45F7BC62") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"30FEF8B580301595353D1056135DD3A6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"85BBEAE208B70D615C45F7BC62";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"30FEF8B580301595353D1056135DD3A6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 459 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"85BBEAE208B70D615C45F7BC62") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8A05B280CA93473356C4290E46BC08AD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"85BBEAE208B70D615C45F7BC62";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8A05B280CA93473356C4290E46BC08AD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 460 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"85BBEAE208B70D615C45F7BC62") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"29BEC9CB33E2844987270ED526887BA8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"85BBEAE208B70D615C45F7BC62";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"29BEC9CB33E2844987270ED526887BA8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 461 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"85BBEAE208B70D615C45F7BC62") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"710FB938DF5D069CF6AD3F0D52420FC3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"85BBEAE208B70D615C45F7BC62";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"710FB938DF5D069CF6AD3F0D52420FC3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 462 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"85BBEAE208B70D615C45F7BC62") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4FC20CAB5577EFF9E60CCB1B0A494F4C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"85BBEAE208B70D615C45F7BC62";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4FC20CAB5577EFF9E60CCB1B0A494F4C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 463 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"85BBEAE208B70D615C45F7BC62D5") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"831EBD7D510E27C22CFC49962F51C7CF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"85BBEAE208B70D615C45F7BC62D5";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"831EBD7D510E27C22CFC49962F51C7CF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 464 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"85BBEAE208B70D615C45F7BC62D5") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5DF03D781CDE54FB11BCA4EFDF767D56") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"85BBEAE208B70D615C45F7BC62D5";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5DF03D781CDE54FB11BCA4EFDF767D56") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 465 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"85BBEAE208B70D615C45F7BC62D5") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7CD8FB56792C185FA80B7DBF5B2E1C89") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"85BBEAE208B70D615C45F7BC62D5";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7CD8FB56792C185FA80B7DBF5B2E1C89") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 466 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"85BBEAE208B70D615C45F7BC62D5") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D84F0AACC1DD252385B904BCAA8FC016") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"85BBEAE208B70D615C45F7BC62D5";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D84F0AACC1DD252385B904BCAA8FC016") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 467 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"85BBEAE208B70D615C45F7BC62D5") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D0C9FB9324C975B1C43E14AB89CBBD25") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"85BBEAE208B70D615C45F7BC62D5";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D0C9FB9324C975B1C43E14AB89CBBD25") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 468 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"85BBEAE208B70D615C45F7BC62D5") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C45AB71F63EC879DBD21EFC361BDE78F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"85BBEAE208B70D615C45F7BC62D5";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C45AB71F63EC879DBD21EFC361BDE78F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 469 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"85BBEAE208B70D615C45F7BC62D5") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F027A6FC1C33E0990F09EAC632F80FDD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"85BBEAE208B70D615C45F7BC62D5";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F027A6FC1C33E0990F09EAC632F80FDD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 470 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"85BBEAE208B70D615C45F7BC62D5") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CDA1D71406F740F9ECCF3831DE70D24D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"85BBEAE208B70D615C45F7BC62D5";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CDA1D71406F740F9ECCF3831DE70D24D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 471 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"85BBEAE208B70D615C45F7BC62D5") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E0533692FC957169E94BDFD33F817783") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"85BBEAE208B70D615C45F7BC62D5";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E0533692FC957169E94BDFD33F817783") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 472 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"85BBEAE208B70D615C45F7BC62D5") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D120F308030A85F14DFF1846392494C3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"85BBEAE208B70D615C45F7BC62D5";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D120F308030A85F14DFF1846392494C3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 473 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"85BBEAE208B70D615C45F7BC62D5") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"22BC92FF118601AFEDBB77161AA2ABCC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"85BBEAE208B70D615C45F7BC62D5";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"22BC92FF118601AFEDBB77161AA2ABCC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 474 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"85BBEAE208B70D615C45F7BC62D5") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"19A079363E7176E90113D9682282F978") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"85BBEAE208B70D615C45F7BC62D5";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"19A079363E7176E90113D9682282F978") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 475 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"85BBEAE208B70D615C45F7BC62D5") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E27136AE313C6B9EDA979F8E87AF2C94") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"85BBEAE208B70D615C45F7BC62D5";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E27136AE313C6B9EDA979F8E87AF2C94") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 476 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"85BBEAE208B70D615C45F7BC62D5") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"681DDF17DBC67BE41C1D93151715790B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"85BBEAE208B70D615C45F7BC62D5";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"681DDF17DBC67BE41C1D93151715790B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 477 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"85BBEAE208B70D615C45F7BC62D5") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"59C78A1FDB773443F48D8CC8C6BEDD8D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"85BBEAE208B70D615C45F7BC62D5";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"59C78A1FDB773443F48D8CC8C6BEDD8D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 478 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"85BBEAE208B70D615C45F7BC62D5") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DC1B5517470CED55F8395743BCFB7A81") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"85BBEAE208B70D615C45F7BC62D5";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DC1B5517470CED55F8395743BCFB7A81") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 479 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"85BBEAE208B70D615C45F7BC62D5") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6C9A0E4AEC0FABD2C01F1625B550325F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"85BBEAE208B70D615C45F7BC62D5";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6C9A0E4AEC0FABD2C01F1625B550325F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 480 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"85BBEAE208B70D615C45F7BC62D5") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D29C369FDFDF69D2386271B78C17B9B5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"85BBEAE208B70D615C45F7BC62D5";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D29C369FDFDF69D2386271B78C17B9B5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 481 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"85BBEAE208B70D615C45F7BC62D5") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"ED32C2F514DF37F99EC5C25ED1B59708") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"85BBEAE208B70D615C45F7BC62D5";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"ED32C2F514DF37F99EC5C25ED1B59708") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 482 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"85BBEAE208B70D615C45F7BC62D5") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7545BADF34CF6C0BE2DBD4800A3BE4D8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"85BBEAE208B70D615C45F7BC62D5";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7545BADF34CF6C0BE2DBD4800A3BE4D8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 483 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"85BBEAE208B70D615C45F7BC62D5") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"09735BEAD071A7A4FFA9C3171448316F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"85BBEAE208B70D615C45F7BC62D5";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"09735BEAD071A7A4FFA9C3171448316F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 484 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"85BBEAE208B70D615C45F7BC62D5") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"09930B31C8D592A0CEB281F49C33F73D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"85BBEAE208B70D615C45F7BC62D5";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"09930B31C8D592A0CEB281F49C33F73D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 485 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"85BBEAE208B70D615C45F7BC62D5") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DA6A9AE77CD3C9D2E4F039E47EBF3FB2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"85BBEAE208B70D615C45F7BC62D5";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DA6A9AE77CD3C9D2E4F039E47EBF3FB2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 486 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"85BBEAE208B70D615C45F7BC62D5") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1C7F9AFD7C9C29B14C6F8F867F230830") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"85BBEAE208B70D615C45F7BC62D5";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1C7F9AFD7C9C29B14C6F8F867F230830") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 487 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"85BBEAE208B70D615C45F7BC62D5") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9A66C211C1EA1FAAAFB5A022583836A6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"85BBEAE208B70D615C45F7BC62D5";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9A66C211C1EA1FAAAFB5A022583836A6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 488 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"85BBEAE208B70D615C45F7BC62D5") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"311D1616C99358D11AF9A82D743490D6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"85BBEAE208B70D615C45F7BC62D5";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"311D1616C99358D11AF9A82D743490D6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 489 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"85BBEAE208B70D615C45F7BC62D5") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"287908E7C8E68301BE63F4570AD3FB96") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"85BBEAE208B70D615C45F7BC62D5";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"287908E7C8E68301BE63F4570AD3FB96") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 490 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"85BBEAE208B70D615C45F7BC62D5") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9DA9F226C632FBC78E068D0B5650DCA5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"85BBEAE208B70D615C45F7BC62D5";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9DA9F226C632FBC78E068D0B5650DCA5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 491 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"85BBEAE208B70D615C45F7BC62D5") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"53D7859C1A766E1988A7E3C77577EFE7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"85BBEAE208B70D615C45F7BC62D5";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"53D7859C1A766E1988A7E3C77577EFE7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 492 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"85BBEAE208B70D615C45F7BC62D5") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E92CCFA950D53CBFEB5EDA9F209634EC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"85BBEAE208B70D615C45F7BC62D5";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E92CCFA950D53CBFEB5EDA9F209634EC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 493 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"85BBEAE208B70D615C45F7BC62D5") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4A97B4E2A9A4FFC53ABDFD4440A247E9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"85BBEAE208B70D615C45F7BC62D5";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4A97B4E2A9A4FFC53ABDFD4440A247E9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 494 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"85BBEAE208B70D615C45F7BC62D5") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1226C411451B7D104B37CC9C34683382") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"85BBEAE208B70D615C45F7BC62D5";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1226C411451B7D104B37CC9C34683382") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 495 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"85BBEAE208B70D615C45F7BC62D5") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2CEB7182CF3194755B96388A6C63730D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"85BBEAE208B70D615C45F7BC62D5";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2CEB7182CF3194755B96388A6C63730D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 496 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"85BBEAE208B70D615C45F7BC62D50D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"38579A311F8B0FB33080A85EE8B61CB6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"85BBEAE208B70D615C45F7BC62D50D";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"38579A311F8B0FB33080A85EE8B61CB6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 497 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"85BBEAE208B70D615C45F7BC62D50D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E6B91A34525B7C8A0DC045271891A62F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"85BBEAE208B70D615C45F7BC62D50D";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E6B91A34525B7C8A0DC045271891A62F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 498 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"85BBEAE208B70D615C45F7BC62D50D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C791DC1A37A9302EB4779C779CC9C7F0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"85BBEAE208B70D615C45F7BC62D50D";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C791DC1A37A9302EB4779C779CC9C7F0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 499 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"85BBEAE208B70D615C45F7BC62D50D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"63062DE08F580D5299C5E5746D681B6F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"85BBEAE208B70D615C45F7BC62D50D";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"63062DE08F580D5299C5E5746D681B6F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      wait;
   end process;

END;
