--
-- SKINNY-AEAD Reference Hardware Implementation
-- 
-- Copyright 2019:
--     Amir Moradi & Pascal Sasdrich for the SKINNY Team
--     https://sites.google.com/site/skinnycipher/
-- 
-- This program is free software; you can redistribute it and/or
-- modify it under the terms of the GNU General Public License as
-- published by the Free Software Foundation; either version 2 of the
-- License, or (at your option) any later version.
-- 
-- This program is distributed in the hope that it will be useful, but
-- WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE. See the GNU
-- General Public License for more details.
-- 

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
ENTITY SKINNY_tk3_AEAD_encdec_M1_Test_Part2 IS
END SKINNY_tk3_AEAD_encdec_M1_Test_Part2;
 
ARCHITECTURE behavior OF SKINNY_tk3_AEAD_encdec_M1_Test_Part2 IS 
 
	constant	nl		 : integer := 0; -- 128-bit nonce
	constant	tl		 : integer := 0; -- 128-bit tag     -> M1
 
 
   COMPONENT SKINNY_tk3_AEAD
	Generic (
		nl				 : integer;  -- 0: 128-bit nonce, 1: 96-bit nonce
		tl				 : integer); -- 0: 128-bit tag,   1: 64-bit tag
	Port (  
		clk          : in  STD_LOGIC;
		rst      	 : in  STD_LOGIC;
		a_data       : in  STD_LOGIC;
		enc          : in  STD_LOGIC;
		dec          : in  STD_LOGIC;
		gen_tag      : in  std_logic;
		Input        : in  STD_LOGIC_VECTOR (127       downto 0);  -- Message or Associated Data
		N            : in  STD_LOGIC_VECTOR (127-nl*32 downto 0);
		K            : in  STD_LOGIC_VECTOR (127       downto 0);
		Block_Size	 : in  STD_LOGIC_VECTOR (  3       downto 0); -- Size of the given block as Input (in BYTES) - 1
		Output       : out STD_LOGIC_VECTOR (127       downto 0); -- Ciphertext
	   Tag			 : out STD_LOGIC_VECTOR (127-tl*64 downto 0); -- Tag
		done         : out STD_LOGIC);
	END COMPONENT;
    

   --Inputs
   signal clk 			: std_logic := '0';
   signal rst 			: std_logic := '0';
   signal a_data 		: std_logic := '0';
   signal enc 			: std_logic := '0';
   signal dec 			: std_logic := '0';
   signal gen_tag 	: std_logic := '0';
   signal Input 		: std_logic_vector(127       downto 0) := (others => '0');
   signal N 			: std_logic_vector(127-nl*32 downto 0) := (others => '0');
   signal K 			: std_logic_vector(127       downto 0) := (others => '0');
   signal Block_Size : std_logic_vector(  3       downto 0) := (others => '0');

 	--Outputs
   signal Output 		: std_logic_vector(127 downto 0);
   signal Tag 		   : std_logic_vector(127-tl*64 downto 0);
   signal done 		: std_logic;

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
   uut: SKINNY_tk3_AEAD 
	GENERIC MAP (
		nl		=> nl,
		tl		=> tl)
	PORT MAP (
		clk 			=> clk,
		rst 			=> rst,
		a_data 		=> a_data,
		enc 			=> enc,
		dec 			=> dec,
		gen_tag 		=> gen_tag,
		Input 		=> Input,
		N 				=> N,
		K 				=> K,
		Block_Size 	=> Block_Size,
		Output 		=> Output,
		Tag			=> Tag,
		done 			=> done);

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      --------- test no. 500 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"85BBEAE208B70D615C45F7BC62D50D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6B80DCDF6A4C5DC0D842F5634E2C665C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"85BBEAE208B70D615C45F7BC62D50D";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6B80DCDF6A4C5DC0D842F5634E2C665C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 501 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"85BBEAE208B70D615C45F7BC62D50D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7F1390532D69AFECA15D0E0BA65A3CF6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"85BBEAE208B70D615C45F7BC62D50D";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7F1390532D69AFECA15D0E0BA65A3CF6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 502 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"85BBEAE208B70D615C45F7BC62D50D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4B6E81B052B6C8E813750B0EF51FD4A4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"85BBEAE208B70D615C45F7BC62D50D";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4B6E81B052B6C8E813750B0EF51FD4A4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 503 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"85BBEAE208B70D615C45F7BC62D50D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"76E8F05848726888F0B3D9F919970934") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"85BBEAE208B70D615C45F7BC62D50D";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"76E8F05848726888F0B3D9F919970934") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 504 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"85BBEAE208B70D615C45F7BC62D50D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5B1A11DEB2105918F5373E1BF866ACFA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"85BBEAE208B70D615C45F7BC62D50D";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5B1A11DEB2105918F5373E1BF866ACFA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 505 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"85BBEAE208B70D615C45F7BC62D50D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6A69D4444D8FAD805183F98EFEC34FBA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"85BBEAE208B70D615C45F7BC62D50D";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6A69D4444D8FAD805183F98EFEC34FBA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 506 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"85BBEAE208B70D615C45F7BC62D50D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"99F5B5B35F0329DEF1C796DEDD4570B5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"85BBEAE208B70D615C45F7BC62D50D";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"99F5B5B35F0329DEF1C796DEDD4570B5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 507 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"85BBEAE208B70D615C45F7BC62D50D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A2E95E7A70F45E981D6F38A0E5652201") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"85BBEAE208B70D615C45F7BC62D50D";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A2E95E7A70F45E981D6F38A0E5652201") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 508 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"85BBEAE208B70D615C45F7BC62D50D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"593811E27FB943EFC6EB7E464048F7ED") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"85BBEAE208B70D615C45F7BC62D50D";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"593811E27FB943EFC6EB7E464048F7ED") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 509 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"85BBEAE208B70D615C45F7BC62D50D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D354F85B95435395006172DDD0F2A272") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"85BBEAE208B70D615C45F7BC62D50D";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D354F85B95435395006172DDD0F2A272") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 510 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"85BBEAE208B70D615C45F7BC62D50D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E28EAD5395F21C32E8F16D00015906F4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"85BBEAE208B70D615C45F7BC62D50D";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E28EAD5395F21C32E8F16D00015906F4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 511 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"85BBEAE208B70D615C45F7BC62D50D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6752725B0989C524E445B68B7B1CA1F8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"85BBEAE208B70D615C45F7BC62D50D";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6752725B0989C524E445B68B7B1CA1F8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 512 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"85BBEAE208B70D615C45F7BC62D50D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D7D32906A28A83A3DC63F7ED72B7E926") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"85BBEAE208B70D615C45F7BC62D50D";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D7D32906A28A83A3DC63F7ED72B7E926") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 513 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"85BBEAE208B70D615C45F7BC62D50D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"69D511D3915A41A3241E907F4BF062CC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"85BBEAE208B70D615C45F7BC62D50D";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"69D511D3915A41A3241E907F4BF062CC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 514 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"85BBEAE208B70D615C45F7BC62D50D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"567BE5B95A5A1F8882B9239616524C71") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"85BBEAE208B70D615C45F7BC62D50D";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"567BE5B95A5A1F8882B9239616524C71") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 515 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"85BBEAE208B70D615C45F7BC62D50D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CE0C9D937A4A447AFEA73548CDDC3FA1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"85BBEAE208B70D615C45F7BC62D50D";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CE0C9D937A4A447AFEA73548CDDC3FA1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 516 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"85BBEAE208B70D615C45F7BC62D50D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B23A7CA69EF48FD5E3D522DFD3AFEA16") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"85BBEAE208B70D615C45F7BC62D50D";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B23A7CA69EF48FD5E3D522DFD3AFEA16") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 517 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"85BBEAE208B70D615C45F7BC62D50D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B2DA2C7D8650BAD1D2CE603C5BD42C44") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"85BBEAE208B70D615C45F7BC62D50D";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B2DA2C7D8650BAD1D2CE603C5BD42C44") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 518 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"85BBEAE208B70D615C45F7BC62D50D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6123BDAB3256E1A3F88CD82CB958E4CB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"85BBEAE208B70D615C45F7BC62D50D";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6123BDAB3256E1A3F88CD82CB958E4CB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 519 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"85BBEAE208B70D615C45F7BC62D50D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A736BDB1321901C050136E4EB8C4D349") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"85BBEAE208B70D615C45F7BC62D50D";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A736BDB1321901C050136E4EB8C4D349") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 520 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"85BBEAE208B70D615C45F7BC62D50D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"212FE55D8F6F37DBB3C941EA9FDFEDDF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"85BBEAE208B70D615C45F7BC62D50D";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"212FE55D8F6F37DBB3C941EA9FDFEDDF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 521 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"85BBEAE208B70D615C45F7BC62D50D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8A54315A871670A0068549E5B3D34BAF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"85BBEAE208B70D615C45F7BC62D50D";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8A54315A871670A0068549E5B3D34BAF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 522 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"85BBEAE208B70D615C45F7BC62D50D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"93302FAB8663AB70A21F159FCD3420EF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"85BBEAE208B70D615C45F7BC62D50D";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"93302FAB8663AB70A21F159FCD3420EF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 523 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"85BBEAE208B70D615C45F7BC62D50D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"26E0D56A88B7D3B6927A6CC391B707DC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"85BBEAE208B70D615C45F7BC62D50D";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"26E0D56A88B7D3B6927A6CC391B707DC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 524 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"85BBEAE208B70D615C45F7BC62D50D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E89EA2D054F3466894DB020FB290349E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"85BBEAE208B70D615C45F7BC62D50D";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E89EA2D054F3466894DB020FB290349E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 525 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"85BBEAE208B70D615C45F7BC62D50D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5265E8E51E5014CEF7223B57E771EF95") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"85BBEAE208B70D615C45F7BC62D50D";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5265E8E51E5014CEF7223B57E771EF95") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 526 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"85BBEAE208B70D615C45F7BC62D50D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F1DE93AEE721D7B426C11C8C87459C90") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"85BBEAE208B70D615C45F7BC62D50D";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F1DE93AEE721D7B426C11C8C87459C90") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 527 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"85BBEAE208B70D615C45F7BC62D50D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A96FE35D0B9E5561574B2D54F38FE8FB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"85BBEAE208B70D615C45F7BC62D50D";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A96FE35D0B9E5561574B2D54F38FE8FB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 528 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"85BBEAE208B70D615C45F7BC62D50D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"97A256CE81B4BC0447EAD942AB84A874") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"85BBEAE208B70D615C45F7BC62D50D";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"97A256CE81B4BC0447EAD942AB84A874") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 529 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B5C35B9E0877404A447206AD8215D411") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B5C35B9E0877404A447206AD8215D411") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 530 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6B2DDB9B45A733737932EBD472326E88") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6B2DDB9B45A733737932EBD472326E88") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 531 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4A051DB520557FD7C0853284F66A0F57") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4A051DB520557FD7C0853284F66A0F57") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 532 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EE92EC4F98A442ABED374B8707CBD3C8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EE92EC4F98A442ABED374B8707CBD3C8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 533 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E6141D707DB01239ACB05B90248FAEFB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E6141D707DB01239ACB05B90248FAEFB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 534 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F28751FC3A95E015D5AFA0F8CCF9F451") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F28751FC3A95E015D5AFA0F8CCF9F451") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 535 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C6FA401F454A87116787A5FD9FBC1C03") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C6FA401F454A87116787A5FD9FBC1C03") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 536 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FB7C31F75F8E27718441770A7334C193") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FB7C31F75F8E27718441770A7334C193") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 537 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D68ED071A5EC16E181C590E892C5645D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D68ED071A5EC16E181C590E892C5645D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 538 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E7FD15EB5A73E2792571577D9460871D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E7FD15EB5A73E2792571577D9460871D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 539 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1461741C48FF66278535382DB7E6B812") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1461741C48FF66278535382DB7E6B812") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 540 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2F7D9FD567081161699D96538FC6EAA6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2F7D9FD567081161699D96538FC6EAA6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 541 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D4ACD04D68450C16B219D0B52AEB3F4A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D4ACD04D68450C16B219D0B52AEB3F4A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 542 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5EC039F482BF1C6C7493DC2EBA516AD5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5EC039F482BF1C6C7493DC2EBA516AD5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 543 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6F1A6CFC820E53CB9C03C3F36BFACE53") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6F1A6CFC820E53CB9C03C3F36BFACE53") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 544 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EAC6B3F41E758ADD90B7187811BF695F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EAC6B3F41E758ADD90B7187811BF695F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 545 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5A47E8A9B576CC5AA891591E18142181") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5A47E8A9B576CC5AA891591E18142181") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 546 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E441D07C86A60E5A50EC3E8C2153AA6B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E441D07C86A60E5A50EC3E8C2153AA6B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 547 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DBEF24164DA65071F64B8D657CF184D6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DBEF24164DA65071F64B8D657CF184D6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 548 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"43985C3C6DB60B838A559BBBA77FF706") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"43985C3C6DB60B838A559BBBA77FF706") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 549 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3FAEBD098908C02C97278C2CB90C22B1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3FAEBD098908C02C97278C2CB90C22B1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 550 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3F4EEDD291ACF528A63CCECF3177E4E3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3F4EEDD291ACF528A63CCECF3177E4E3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 551 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"ECB77C0425AAAE5A8C7E76DFD3FB2C6C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"ECB77C0425AAAE5A8C7E76DFD3FB2C6C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 552 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2AA27C1E25E54E3924E1C0BDD2671BEE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2AA27C1E25E54E3924E1C0BDD2671BEE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 553 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"ACBB24F298937822C73BEF19F57C2578") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"ACBB24F298937822C73BEF19F57C2578") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 554 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"07C0F0F590EA3F597277E716D9708308") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"07C0F0F590EA3F597277E716D9708308") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 555 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1EA4EE04919FE489D6EDBB6CA797E848") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1EA4EE04919FE489D6EDBB6CA797E848") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 556 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AB7414C59F4B9C4FE688C230FB14CF7B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AB7414C59F4B9C4FE688C230FB14CF7B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 557 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"650A637F430F0991E029ACFCD833FC39") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"650A637F430F0991E029ACFCD833FC39") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 558 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DFF1294A09AC5B3783D095A48DD22732") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DFF1294A09AC5B3783D095A48DD22732") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 559 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7C4A5201F0DD984D5233B27FEDE65437") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7C4A5201F0DD984D5233B27FEDE65437") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 560 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"24FB22F21C621A9823B983A7992C205C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"24FB22F21C621A9823B983A7992C205C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 561 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1A3697619648F3FD331877B1C12760D3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1A3697619648F3FD331877B1C12760D3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 562 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"9A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AFFCC7BE1FD1B7101D287E7179FA49B5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"9A";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AFFCC7BE1FD1B7101D287E7179FA49B5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 563 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"9A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"711247BB5201C4292068930889DDF32C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"9A";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"711247BB5201C4292068930889DDF32C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 564 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"9A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"503A819537F3888D99DF4A580D8592F3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"9A";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"503A819537F3888D99DF4A580D8592F3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 565 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"9A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F4AD706F8F02B5F1B46D335BFC244E6C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"9A";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F4AD706F8F02B5F1B46D335BFC244E6C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 566 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"9A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FC2B81506A16E563F5EA234CDF60335F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"9A";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FC2B81506A16E563F5EA234CDF60335F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 567 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"9A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E8B8CDDC2D33174F8CF5D824371669F5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"9A";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E8B8CDDC2D33174F8CF5D824371669F5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 568 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"9A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DCC5DC3F52EC704B3EDDDD21645381A7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"9A";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DCC5DC3F52EC704B3EDDDD21645381A7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 569 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"9A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E143ADD74828D02BDD1B0FD688DB5C37") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"9A";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E143ADD74828D02BDD1B0FD688DB5C37") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 570 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"9A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CCB14C51B24AE1BBD89FE834692AF9F9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"9A";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CCB14C51B24AE1BBD89FE834692AF9F9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 571 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"9A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FDC289CB4DD515237C2B2FA16F8F1AB9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"9A";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FDC289CB4DD515237C2B2FA16F8F1AB9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 572 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"9A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0E5EE83C5F59917DDC6F40F14C0925B6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"9A";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0E5EE83C5F59917DDC6F40F14C0925B6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 573 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"9A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"354203F570AEE63B30C7EE8F74297702") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"9A";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"354203F570AEE63B30C7EE8F74297702") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 574 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"9A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CE934C6D7FE3FB4CEB43A869D104A2EE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"9A";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CE934C6D7FE3FB4CEB43A869D104A2EE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 575 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"9A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"44FFA5D49519EB362DC9A4F241BEF771") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"9A";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"44FFA5D49519EB362DC9A4F241BEF771") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 576 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"9A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7525F0DC95A8A491C559BB2F901553F7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"9A";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7525F0DC95A8A491C559BB2F901553F7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 577 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"9A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F0F92FD409D37D87C9ED60A4EA50F4FB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"9A";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F0F92FD409D37D87C9ED60A4EA50F4FB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 578 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"9A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"40787489A2D03B00F1CB21C2E3FBBC25") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"9A";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"40787489A2D03B00F1CB21C2E3FBBC25") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 579 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"9A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FE7E4C5C9100F90009B64650DABC37CF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"9A";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FE7E4C5C9100F90009B64650DABC37CF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 580 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"9A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C1D0B8365A00A72BAF11F5B9871E1972") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"9A";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C1D0B8365A00A72BAF11F5B9871E1972") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 581 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"9A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"59A7C01C7A10FCD9D30FE3675C906AA2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"9A";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"59A7C01C7A10FCD9D30FE3675C906AA2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 582 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"9A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"259121299EAE3776CE7DF4F042E3BF15") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"9A";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"259121299EAE3776CE7DF4F042E3BF15") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 583 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"9A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"257171F2860A0272FF66B613CA987947") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"9A";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"257171F2860A0272FF66B613CA987947") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 584 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"9A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F688E024320C5900D5240E032814B1C8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"9A";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F688E024320C5900D5240E032814B1C8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 585 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"9A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"309DE03E3243B9637DBBB8612988864A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"9A";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"309DE03E3243B9637DBBB8612988864A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 586 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"9A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B684B8D28F358F789E6197C50E93B8DC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"9A";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B684B8D28F358F789E6197C50E93B8DC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 587 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"9A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1DFF6CD5874CC8032B2D9FCA229F1EAC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"9A";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1DFF6CD5874CC8032B2D9FCA229F1EAC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 588 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"9A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"049B7224863913D38FB7C3B05C7875EC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"9A";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"049B7224863913D38FB7C3B05C7875EC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 589 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"9A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B14B88E588ED6B15BFD2BAEC00FB52DF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"9A";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B14B88E588ED6B15BFD2BAEC00FB52DF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 590 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"9A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7F35FF5F54A9FECBB973D42023DC619D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"9A";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7F35FF5F54A9FECBB973D42023DC619D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 591 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"9A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C5CEB56A1E0AAC6DDA8AED78763DBA96") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"9A";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C5CEB56A1E0AAC6DDA8AED78763DBA96") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 592 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"9A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6675CE21E77B6F170B69CAA31609C993") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"9A";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6675CE21E77B6F170B69CAA31609C993") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 593 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"9A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3EC4BED20BC4EDC27AE3FB7B62C3BDF8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"9A";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3EC4BED20BC4EDC27AE3FB7B62C3BDF8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 594 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"9A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"00090B4181EE04A76A420F6D3AC8FD77") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"9A";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"00090B4181EE04A76A420F6D3AC8FD77") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 595 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"9A15") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BCD31E9BCE28BE30DD35DC07BFE893DF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"9A15";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BCD31E9BCE28BE30DD35DC07BFE893DF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 596 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"9A15") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"623D9E9E83F8CD09E075317E4FCF2946") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"9A15";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"623D9E9E83F8CD09E075317E4FCF2946") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 597 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"9A15") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"431558B0E60A81AD59C2E82ECB974899") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"9A15";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"431558B0E60A81AD59C2E82ECB974899") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 598 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"9A15") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E782A94A5EFBBCD17470912D3A369406") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"9A15";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E782A94A5EFBBCD17470912D3A369406") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 599 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"9A15") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EF045875BBEFEC4335F7813A1972E935") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"9A15";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EF045875BBEFEC4335F7813A1972E935") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 600 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"9A15") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FB9714F9FCCA1E6F4CE87A52F104B39F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"9A15";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FB9714F9FCCA1E6F4CE87A52F104B39F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 601 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"9A15") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CFEA051A8315796BFEC07F57A2415BCD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"9A15";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CFEA051A8315796BFEC07F57A2415BCD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 602 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"9A15") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F26C74F299D1D90B1D06ADA04EC9865D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"9A15";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F26C74F299D1D90B1D06ADA04EC9865D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 603 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"9A15") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DF9E957463B3E89B18824A42AF382393") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"9A15";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DF9E957463B3E89B18824A42AF382393") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 604 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"9A15") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EEED50EE9C2C1C03BC368DD7A99DC0D3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"9A15";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EEED50EE9C2C1C03BC368DD7A99DC0D3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 605 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"9A15") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1D7131198EA0985D1C72E2878A1BFFDC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"9A15";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1D7131198EA0985D1C72E2878A1BFFDC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 606 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"9A15") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"266DDAD0A157EF1BF0DA4CF9B23BAD68") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"9A15";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"266DDAD0A157EF1BF0DA4CF9B23BAD68") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 607 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"9A15") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DDBC9548AE1AF26C2B5E0A1F17167884") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"9A15";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DDBC9548AE1AF26C2B5E0A1F17167884") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 608 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"9A15") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"57D07CF144E0E216EDD4068487AC2D1B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"9A15";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"57D07CF144E0E216EDD4068487AC2D1B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 609 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"9A15") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"660A29F94451ADB1054419595607899D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"9A15";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"660A29F94451ADB1054419595607899D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 610 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"9A15") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E3D6F6F1D82A74A709F0C2D22C422E91") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"9A15";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E3D6F6F1D82A74A709F0C2D22C422E91") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 611 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"9A15") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5357ADAC7329322031D683B425E9664F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"9A15";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5357ADAC7329322031D683B425E9664F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 612 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"9A15") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"ED51957940F9F020C9ABE4261CAEEDA5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"9A15";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"ED51957940F9F020C9ABE4261CAEEDA5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 613 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"9A15") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D2FF61138BF9AE0B6F0C57CF410CC318") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"9A15";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D2FF61138BF9AE0B6F0C57CF410CC318") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 614 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"9A15") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4A881939ABE9F5F9131241119A82B0C8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"9A15";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4A881939ABE9F5F9131241119A82B0C8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 615 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"9A15") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"36BEF80C4F573E560E60568684F1657F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"9A15";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"36BEF80C4F573E560E60568684F1657F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 616 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"9A15") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"365EA8D757F30B523F7B14650C8AA32D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"9A15";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"365EA8D757F30B523F7B14650C8AA32D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 617 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"9A15") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E5A73901E3F550201539AC75EE066BA2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"9A15";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E5A73901E3F550201539AC75EE066BA2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 618 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"9A15") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"23B2391BE3BAB043BDA61A17EF9A5C20") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"9A15";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"23B2391BE3BAB043BDA61A17EF9A5C20") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 619 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"9A15") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A5AB61F75ECC86585E7C35B3C88162B6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"9A15";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A5AB61F75ECC86585E7C35B3C88162B6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 620 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"9A15") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0ED0B5F056B5C123EB303DBCE48DC4C6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"9A15";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0ED0B5F056B5C123EB303DBCE48DC4C6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 621 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"9A15") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"17B4AB0157C01AF34FAA61C69A6AAF86") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"9A15";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"17B4AB0157C01AF34FAA61C69A6AAF86") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 622 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"9A15") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A26451C0591462357FCF189AC6E988B5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"9A15";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A26451C0591462357FCF189AC6E988B5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 623 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"9A15") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6C1A267A8550F7EB796E7656E5CEBBF7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"9A15";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6C1A267A8550F7EB796E7656E5CEBBF7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 624 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"9A15") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D6E16C4FCFF3A54D1A974F0EB02F60FC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"9A15";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D6E16C4FCFF3A54D1A974F0EB02F60FC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 625 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"9A15") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"755A170436826637CB7468D5D01B13F9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"9A15";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"755A170436826637CB7468D5D01B13F9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 626 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"9A15") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2DEB67F7DA3DE4E2BAFE590DA4D16792") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"9A15";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2DEB67F7DA3DE4E2BAFE590DA4D16792") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 627 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"9A15") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1326D26450170D87AA5FAD1BFCDA271D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"9A15";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1326D26450170D87AA5FAD1BFCDA271D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 628 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"9A1562") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3FDADA47D472EE1907F501BEBA07366E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"9A1562";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3FDADA47D472EE1907F501BEBA07366E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 629 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"9A1562") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E1345A4299A29D203AB5ECC74A208CF7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"9A1562";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E1345A4299A29D203AB5ECC74A208CF7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 630 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"9A1562") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C01C9C6CFC50D18483023597CE78ED28") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"9A1562";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C01C9C6CFC50D18483023597CE78ED28") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 631 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"9A1562") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"648B6D9644A1ECF8AEB04C943FD931B7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"9A1562";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"648B6D9644A1ECF8AEB04C943FD931B7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 632 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"9A1562") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6C0D9CA9A1B5BC6AEF375C831C9D4C84") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"9A1562";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6C0D9CA9A1B5BC6AEF375C831C9D4C84") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 633 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"9A1562") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"789ED025E6904E469628A7EBF4EB162E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"9A1562";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"789ED025E6904E469628A7EBF4EB162E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 634 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"9A1562") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4CE3C1C6994F29422400A2EEA7AEFE7C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"9A1562";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4CE3C1C6994F29422400A2EEA7AEFE7C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 635 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"9A1562") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7165B02E838B8922C7C670194B2623EC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"9A1562";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7165B02E838B8922C7C670194B2623EC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 636 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"9A1562") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5C9751A879E9B8B2C24297FBAAD78622") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"9A1562";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5C9751A879E9B8B2C24297FBAAD78622") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 637 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"9A1562") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6DE4943286764C2A66F6506EAC726562") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"9A1562";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6DE4943286764C2A66F6506EAC726562") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 638 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"9A1562") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9E78F5C594FAC874C6B23F3E8FF45A6D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"9A1562";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9E78F5C594FAC874C6B23F3E8FF45A6D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 639 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"9A1562") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A5641E0CBB0DBF322A1A9140B7D408D9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"9A1562";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A5641E0CBB0DBF322A1A9140B7D408D9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 640 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"9A1562") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5EB55194B440A245F19ED7A612F9DD35") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"9A1562";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5EB55194B440A245F19ED7A612F9DD35") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 641 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"9A1562") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D4D9B82D5EBAB23F3714DB3D824388AA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"9A1562";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D4D9B82D5EBAB23F3714DB3D824388AA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 642 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"9A1562") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E503ED255E0BFD98DF84C4E053E82C2C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"9A1562";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E503ED255E0BFD98DF84C4E053E82C2C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 643 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"9A1562") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"60DF322DC270248ED3301F6B29AD8B20") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"9A1562";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"60DF322DC270248ED3301F6B29AD8B20") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 644 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"9A1562") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D05E697069736209EB165E0D2006C3FE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"9A1562";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D05E697069736209EB165E0D2006C3FE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 645 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"9A1562") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6E5851A55AA3A009136B399F19414814") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"9A1562";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6E5851A55AA3A009136B399F19414814") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 646 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"9A1562") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"51F6A5CF91A3FE22B5CC8A7644E366A9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"9A1562";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"51F6A5CF91A3FE22B5CC8A7644E366A9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 647 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"9A1562") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C981DDE5B1B3A5D0C9D29CA89F6D1579") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"9A1562";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C981DDE5B1B3A5D0C9D29CA89F6D1579") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 648 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"9A1562") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B5B73CD0550D6E7FD4A08B3F811EC0CE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"9A1562";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B5B73CD0550D6E7FD4A08B3F811EC0CE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 649 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"9A1562") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B5576C0B4DA95B7BE5BBC9DC0965069C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"9A1562";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B5576C0B4DA95B7BE5BBC9DC0965069C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 650 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"9A1562") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"66AEFDDDF9AF0009CFF971CCEBE9CE13") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"9A1562";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"66AEFDDDF9AF0009CFF971CCEBE9CE13") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 651 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"9A1562") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A0BBFDC7F9E0E06A6766C7AEEA75F991") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"9A1562";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A0BBFDC7F9E0E06A6766C7AEEA75F991") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 652 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"9A1562") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"26A2A52B4496D67184BCE80ACD6EC707") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"9A1562";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"26A2A52B4496D67184BCE80ACD6EC707") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 653 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"9A1562") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8DD9712C4CEF910A31F0E005E1626177") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"9A1562";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8DD9712C4CEF910A31F0E005E1626177") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 654 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"9A1562") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"94BD6FDD4D9A4ADA956ABC7F9F850A37") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"9A1562";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"94BD6FDD4D9A4ADA956ABC7F9F850A37") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 655 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"9A1562") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"216D951C434E321CA50FC523C3062D04") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"9A1562";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"216D951C434E321CA50FC523C3062D04") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 656 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"9A1562") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EF13E2A69F0AA7C2A3AEABEFE0211E46") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"9A1562";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EF13E2A69F0AA7C2A3AEABEFE0211E46") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 657 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"9A1562") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"55E8A893D5A9F564C05792B7B5C0C54D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"9A1562";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"55E8A893D5A9F564C05792B7B5C0C54D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 658 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"9A1562") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F653D3D82CD8361E11B4B56CD5F4B648") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"9A1562";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F653D3D82CD8361E11B4B56CD5F4B648") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 659 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"9A1562") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AEE2A32BC067B4CB603E84B4A13EC223") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"9A1562";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AEE2A32BC067B4CB603E84B4A13EC223") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 660 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"9A1562") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"902F16B84A4D5DAE709F70A2F93582AC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"9A1562";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"902F16B84A4D5DAE709F70A2F93582AC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 661 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"9A1562B4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FF116C4E5E99F61BA9F5EDD799EB4D44") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"9A1562B4";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FF116C4E5E99F61BA9F5EDD799EB4D44") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 662 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"9A1562B4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"21FFEC4B1349852294B500AE69CCF7DD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"9A1562B4";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"21FFEC4B1349852294B500AE69CCF7DD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 663 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"9A1562B4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"00D72A6576BBC9862D02D9FEED949602") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"9A1562B4";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"00D72A6576BBC9862D02D9FEED949602") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 664 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"9A1562B4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A440DB9FCE4AF4FA00B0A0FD1C354A9D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"9A1562B4";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A440DB9FCE4AF4FA00B0A0FD1C354A9D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 665 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"9A1562B4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"ACC62AA02B5EA4684137B0EA3F7137AE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"9A1562B4";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"ACC62AA02B5EA4684137B0EA3F7137AE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 666 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"9A1562B4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B855662C6C7B564438284B82D7076D04") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"9A1562B4";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B855662C6C7B564438284B82D7076D04") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 667 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"9A1562B4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8C2877CF13A431408A004E8784428556") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"9A1562B4";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8C2877CF13A431408A004E8784428556") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 668 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"9A1562B4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B1AE06270960912069C69C7068CA58C6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"9A1562B4";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B1AE06270960912069C69C7068CA58C6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 669 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"9A1562B4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9C5CE7A1F302A0B06C427B92893BFD08") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"9A1562B4";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9C5CE7A1F302A0B06C427B92893BFD08") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 670 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"9A1562B4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AD2F223B0C9D5428C8F6BC078F9E1E48") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"9A1562B4";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AD2F223B0C9D5428C8F6BC078F9E1E48") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 671 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"9A1562B4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5EB343CC1E11D07668B2D357AC182147") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"9A1562B4";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5EB343CC1E11D07668B2D357AC182147") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 672 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"9A1562B4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"65AFA80531E6A730841A7D29943873F3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"9A1562B4";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"65AFA80531E6A730841A7D29943873F3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 673 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"9A1562B4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9E7EE79D3EABBA475F9E3BCF3115A61F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"9A1562B4";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9E7EE79D3EABBA475F9E3BCF3115A61F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 674 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"9A1562B4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"14120E24D451AA3D99143754A1AFF380") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"9A1562B4";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"14120E24D451AA3D99143754A1AFF380") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 675 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"9A1562B4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"25C85B2CD4E0E59A7184288970045706") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"9A1562B4";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"25C85B2CD4E0E59A7184288970045706") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 676 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"9A1562B4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A0148424489B3C8C7D30F3020A41F00A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"9A1562B4";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A0148424489B3C8C7D30F3020A41F00A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 677 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"9A1562B4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1095DF79E3987A0B4516B26403EAB8D4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"9A1562B4";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1095DF79E3987A0B4516B26403EAB8D4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 678 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"9A1562B4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AE93E7ACD048B80BBD6BD5F63AAD333E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"9A1562B4";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AE93E7ACD048B80BBD6BD5F63AAD333E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 679 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"9A1562B4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"913D13C61B48E6201BCC661F670F1D83") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"9A1562B4";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"913D13C61B48E6201BCC661F670F1D83") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 680 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"9A1562B4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"094A6BEC3B58BDD267D270C1BC816E53") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"9A1562B4";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"094A6BEC3B58BDD267D270C1BC816E53") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 681 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"9A1562B4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"757C8AD9DFE6767D7AA06756A2F2BBE4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"9A1562B4";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"757C8AD9DFE6767D7AA06756A2F2BBE4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 682 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"9A1562B4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"759CDA02C74243794BBB25B52A897DB6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"9A1562B4";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"759CDA02C74243794BBB25B52A897DB6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 683 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"9A1562B4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A6654BD47344180B61F99DA5C805B539") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"9A1562B4";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A6654BD47344180B61F99DA5C805B539") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 684 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"9A1562B4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"60704BCE730BF868C9662BC7C99982BB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"9A1562B4";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"60704BCE730BF868C9662BC7C99982BB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 685 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"9A1562B4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E6691322CE7DCE732ABC0463EE82BC2D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"9A1562B4";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E6691322CE7DCE732ABC0463EE82BC2D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 686 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"9A1562B4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4D12C725C60489089FF00C6CC28E1A5D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"9A1562B4";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4D12C725C60489089FF00C6CC28E1A5D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 687 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"9A1562B4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5476D9D4C77152D83B6A5016BC69711D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"9A1562B4";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5476D9D4C77152D83B6A5016BC69711D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 688 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"9A1562B4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E1A62315C9A52A1E0B0F294AE0EA562E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"9A1562B4";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E1A62315C9A52A1E0B0F294AE0EA562E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 689 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"9A1562B4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2FD854AF15E1BFC00DAE4786C3CD656C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"9A1562B4";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2FD854AF15E1BFC00DAE4786C3CD656C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 690 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"9A1562B4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"95231E9A5F42ED666E577EDE962CBE67") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"9A1562B4";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"95231E9A5F42ED666E577EDE962CBE67") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 691 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"9A1562B4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"369865D1A6332E1CBFB45905F618CD62") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"9A1562B4";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"369865D1A6332E1CBFB45905F618CD62") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 692 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"9A1562B4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6E2915224A8CACC9CE3E68DD82D2B909") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"9A1562B4";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6E2915224A8CACC9CE3E68DD82D2B909") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 693 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"9A1562B4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"50E4A0B1C0A645ACDE9F9CCBDAD9F986") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"9A1562B4";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"50E4A0B1C0A645ACDE9F9CCBDAD9F986") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 694 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"9A1562B41D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6619BF751B84E0CC84D3CF93160199AD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"9A1562B41D";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6619BF751B84E0CC84D3CF93160199AD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 695 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"9A1562B41D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B8F73F70565493F5B99322EAE6262334") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"9A1562B41D";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B8F73F70565493F5B99322EAE6262334") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 696 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"9A1562B41D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"99DFF95E33A6DF510024FBBA627E42EB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"9A1562B41D";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"99DFF95E33A6DF510024FBBA627E42EB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 697 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"9A1562B41D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3D4808A48B57E22D2D9682B993DF9E74") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"9A1562B41D";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3D4808A48B57E22D2D9682B993DF9E74") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 698 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"9A1562B41D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"35CEF99B6E43B2BF6C1192AEB09BE347") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"9A1562B41D";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"35CEF99B6E43B2BF6C1192AEB09BE347") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 699 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"9A1562B41D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"215DB51729664093150E69C658EDB9ED") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"9A1562B41D";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"215DB51729664093150E69C658EDB9ED") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 700 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"9A1562B41D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1520A4F456B92797A7266CC30BA851BF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"9A1562B41D";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1520A4F456B92797A7266CC30BA851BF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 701 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"9A1562B41D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"28A6D51C4C7D87F744E0BE34E7208C2F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"9A1562B41D";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"28A6D51C4C7D87F744E0BE34E7208C2F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 702 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"9A1562B41D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0554349AB61FB667416459D606D129E1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"9A1562B41D";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0554349AB61FB667416459D606D129E1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 703 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"9A1562B41D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3427F100498042FFE5D09E430074CAA1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"9A1562B41D";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3427F100498042FFE5D09E430074CAA1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 704 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"9A1562B41D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C7BB90F75B0CC6A14594F11323F2F5AE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"9A1562B41D";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C7BB90F75B0CC6A14594F11323F2F5AE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 705 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"9A1562B41D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FCA77B3E74FBB1E7A93C5F6D1BD2A71A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"9A1562B41D";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FCA77B3E74FBB1E7A93C5F6D1BD2A71A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 706 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"9A1562B41D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"077634A67BB6AC9072B8198BBEFF72F6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"9A1562B41D";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"077634A67BB6AC9072B8198BBEFF72F6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 707 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"9A1562B41D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8D1ADD1F914CBCEAB43215102E452769") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"9A1562B41D";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8D1ADD1F914CBCEAB43215102E452769") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 708 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"9A1562B41D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BCC0881791FDF34D5CA20ACDFFEE83EF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"9A1562B41D";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BCC0881791FDF34D5CA20ACDFFEE83EF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 709 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"9A1562B41D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"391C571F0D862A5B5016D14685AB24E3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"9A1562B41D";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"391C571F0D862A5B5016D14685AB24E3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 710 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"9A1562B41D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"899D0C42A6856CDC683090208C006C3D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"9A1562B41D";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"899D0C42A6856CDC683090208C006C3D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 711 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"9A1562B41D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"379B34979555AEDC904DF7B2B547E7D7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"9A1562B41D";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"379B34979555AEDC904DF7B2B547E7D7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 712 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"9A1562B41D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0835C0FD5E55F0F736EA445BE8E5C96A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"9A1562B41D";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0835C0FD5E55F0F736EA445BE8E5C96A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 713 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"9A1562B41D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9042B8D77E45AB054AF45285336BBABA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"9A1562B41D";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9042B8D77E45AB054AF45285336BBABA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 714 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"9A1562B41D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EC7459E29AFB60AA578645122D186F0D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"9A1562B41D";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EC7459E29AFB60AA578645122D186F0D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 715 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"9A1562B41D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EC940939825F55AE669D07F1A563A95F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"9A1562B41D";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EC940939825F55AE669D07F1A563A95F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 716 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"9A1562B41D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3F6D98EF36590EDC4CDFBFE147EF61D0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"9A1562B41D";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3F6D98EF36590EDC4CDFBFE147EF61D0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 717 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"9A1562B41D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F97898F53616EEBFE440098346735652") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"9A1562B41D";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F97898F53616EEBFE440098346735652") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 718 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"9A1562B41D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7F61C0198B60D8A4079A2627616868C4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"9A1562B41D";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7F61C0198B60D8A4079A2627616868C4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 719 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"9A1562B41D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D41A141E83199FDFB2D62E284D64CEB4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"9A1562B41D";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D41A141E83199FDFB2D62E284D64CEB4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 720 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"9A1562B41D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CD7E0AEF826C440F164C72523383A5F4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"9A1562B41D";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CD7E0AEF826C440F164C72523383A5F4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 721 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"9A1562B41D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"78AEF02E8CB83CC926290B0E6F0082C7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"9A1562B41D";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"78AEF02E8CB83CC926290B0E6F0082C7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 722 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"9A1562B41D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B6D0879450FCA917208865C24C27B185") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"9A1562B41D";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B6D0879450FCA917208865C24C27B185") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 723 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"9A1562B41D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0C2BCDA11A5FFBB143715C9A19C66A8E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"9A1562B41D";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0C2BCDA11A5FFBB143715C9A19C66A8E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 724 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"9A1562B41D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AF90B6EAE32E38CB92927B4179F2198B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"9A1562B41D";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AF90B6EAE32E38CB92927B4179F2198B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 725 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"9A1562B41D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F721C6190F91BA1EE3184A990D386DE0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"9A1562B41D";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F721C6190F91BA1EE3184A990D386DE0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 726 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"9A1562B41D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C9EC738A85BB537BF3B9BE8F55332D6F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"9A1562B41D";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C9EC738A85BB537BF3B9BE8F55332D6F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 727 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"9A1562B41DFC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"78A4DF18B1A8D0DD9A93B16EEE3FAD4E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"9A1562B41DFC";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"78A4DF18B1A8D0DD9A93B16EEE3FAD4E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 728 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"9A1562B41DFC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A64A5F1DFC78A3E4A7D35C171E1817D7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"9A1562B41DFC";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A64A5F1DFC78A3E4A7D35C171E1817D7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 729 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"9A1562B41DFC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"87629933998AEF401E6485479A407608") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"9A1562B41DFC";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"87629933998AEF401E6485479A407608") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 730 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"9A1562B41DFC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"23F568C9217BD23C33D6FC446BE1AA97") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"9A1562B41DFC";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"23F568C9217BD23C33D6FC446BE1AA97") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 731 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"9A1562B41DFC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2B7399F6C46F82AE7251EC5348A5D7A4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"9A1562B41DFC";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2B7399F6C46F82AE7251EC5348A5D7A4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 732 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"9A1562B41DFC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3FE0D57A834A70820B4E173BA0D38D0E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"9A1562B41DFC";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3FE0D57A834A70820B4E173BA0D38D0E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 733 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"9A1562B41DFC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0B9DC499FC951786B966123EF396655C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"9A1562B41DFC";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0B9DC499FC951786B966123EF396655C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 734 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"9A1562B41DFC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"361BB571E651B7E65AA0C0C91F1EB8CC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"9A1562B41DFC";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"361BB571E651B7E65AA0C0C91F1EB8CC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 735 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"9A1562B41DFC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1BE954F71C3386765F24272BFEEF1D02") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"9A1562B41DFC";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1BE954F71C3386765F24272BFEEF1D02") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 736 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"9A1562B41DFC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2A9A916DE3AC72EEFB90E0BEF84AFE42") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"9A1562B41DFC";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2A9A916DE3AC72EEFB90E0BEF84AFE42") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 737 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"9A1562B41DFC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D906F09AF120F6B05BD48FEEDBCCC14D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"9A1562B41DFC";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D906F09AF120F6B05BD48FEEDBCCC14D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 738 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"9A1562B41DFC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E21A1B53DED781F6B77C2190E3EC93F9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"9A1562B41DFC";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E21A1B53DED781F6B77C2190E3EC93F9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 739 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"9A1562B41DFC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"19CB54CBD19A9C816CF8677646C14615") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"9A1562B41DFC";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"19CB54CBD19A9C816CF8677646C14615") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 740 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"9A1562B41DFC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"93A7BD723B608CFBAA726BEDD67B138A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"9A1562B41DFC";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"93A7BD723B608CFBAA726BEDD67B138A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 741 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"9A1562B41DFC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A27DE87A3BD1C35C42E2743007D0B70C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"9A1562B41DFC";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A27DE87A3BD1C35C42E2743007D0B70C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 742 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"9A1562B41DFC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"27A13772A7AA1A4A4E56AFBB7D951000") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"9A1562B41DFC";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"27A13772A7AA1A4A4E56AFBB7D951000") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 743 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"9A1562B41DFC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"97206C2F0CA95CCD7670EEDD743E58DE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"9A1562B41DFC";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"97206C2F0CA95CCD7670EEDD743E58DE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 744 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"9A1562B41DFC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"292654FA3F799ECD8E0D894F4D79D334") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"9A1562B41DFC";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"292654FA3F799ECD8E0D894F4D79D334") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 745 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"9A1562B41DFC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1688A090F479C0E628AA3AA610DBFD89") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"9A1562B41DFC";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1688A090F479C0E628AA3AA610DBFD89") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 746 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"9A1562B41DFC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8EFFD8BAD4699B1454B42C78CB558E59") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"9A1562B41DFC";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8EFFD8BAD4699B1454B42C78CB558E59") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 747 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"9A1562B41DFC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F2C9398F30D750BB49C63BEFD5265BEE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"9A1562B41DFC";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F2C9398F30D750BB49C63BEFD5265BEE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 748 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"9A1562B41DFC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F2296954287365BF78DD790C5D5D9DBC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"9A1562B41DFC";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F2296954287365BF78DD790C5D5D9DBC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 749 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"9A1562B41DFC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"21D0F8829C753ECD529FC11CBFD15533") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"9A1562B41DFC";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"21D0F8829C753ECD529FC11CBFD15533") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 750 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"9A1562B41DFC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E7C5F8989C3ADEAEFA00777EBE4D62B1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"9A1562B41DFC";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E7C5F8989C3ADEAEFA00777EBE4D62B1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 751 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"9A1562B41DFC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"61DCA074214CE8B519DA58DA99565C27") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"9A1562B41DFC";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"61DCA074214CE8B519DA58DA99565C27") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 752 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"9A1562B41DFC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CAA774732935AFCEAC9650D5B55AFA57") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"9A1562B41DFC";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CAA774732935AFCEAC9650D5B55AFA57") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 753 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"9A1562B41DFC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D3C36A822840741E080C0CAFCBBD9117") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"9A1562B41DFC";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D3C36A822840741E080C0CAFCBBD9117") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 754 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"9A1562B41DFC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6613904326940CD8386975F3973EB624") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"9A1562B41DFC";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6613904326940CD8386975F3973EB624") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 755 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"9A1562B41DFC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A86DE7F9FAD099063EC81B3FB4198566") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"9A1562B41DFC";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A86DE7F9FAD099063EC81B3FB4198566") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 756 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"9A1562B41DFC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1296ADCCB073CBA05D312267E1F85E6D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"9A1562B41DFC";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1296ADCCB073CBA05D312267E1F85E6D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 757 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"9A1562B41DFC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B12DD687490208DA8CD205BC81CC2D68") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"9A1562B41DFC";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B12DD687490208DA8CD205BC81CC2D68") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 758 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"9A1562B41DFC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E99CA674A5BD8A0FFD583464F5065903") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"9A1562B41DFC";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E99CA674A5BD8A0FFD583464F5065903") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 759 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"9A1562B41DFC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D75113E72F97636AEDF9C072AD0D198C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"9A1562B41DFC";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D75113E72F97636AEDF9C072AD0D198C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 760 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"9A1562B41DFC09") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6DBAC73BCBBB2875C88FFABA25C3FF8B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"9A1562B41DFC09";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6DBAC73BCBBB2875C88FFABA25C3FF8B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 761 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"9A1562B41DFC09") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B354473E866B5B4CF5CF17C3D5E44512") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"9A1562B41DFC09";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B354473E866B5B4CF5CF17C3D5E44512") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 762 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"9A1562B41DFC09") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"927C8110E39917E84C78CE9351BC24CD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"9A1562B41DFC09";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"927C8110E39917E84C78CE9351BC24CD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 763 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"9A1562B41DFC09") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"36EB70EA5B682A9461CAB790A01DF852") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"9A1562B41DFC09";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"36EB70EA5B682A9461CAB790A01DF852") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 764 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"9A1562B41DFC09") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3E6D81D5BE7C7A06204DA78783598561") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"9A1562B41DFC09";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3E6D81D5BE7C7A06204DA78783598561") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 765 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"9A1562B41DFC09") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2AFECD59F959882A59525CEF6B2FDFCB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"9A1562B41DFC09";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2AFECD59F959882A59525CEF6B2FDFCB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 766 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"9A1562B41DFC09") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1E83DCBA8686EF2EEB7A59EA386A3799") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"9A1562B41DFC09";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1E83DCBA8686EF2EEB7A59EA386A3799") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 767 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"9A1562B41DFC09") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2305AD529C424F4E08BC8B1DD4E2EA09") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"9A1562B41DFC09";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2305AD529C424F4E08BC8B1DD4E2EA09") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 768 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"9A1562B41DFC09") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0EF74CD466207EDE0D386CFF35134FC7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"9A1562B41DFC09";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0EF74CD466207EDE0D386CFF35134FC7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 769 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"9A1562B41DFC09") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3F84894E99BF8A46A98CAB6A33B6AC87") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"9A1562B41DFC09";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3F84894E99BF8A46A98CAB6A33B6AC87") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 770 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"9A1562B41DFC09") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CC18E8B98B330E1809C8C43A10309388") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"9A1562B41DFC09";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CC18E8B98B330E1809C8C43A10309388") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 771 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"9A1562B41DFC09") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F7040370A4C4795EE5606A442810C13C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"9A1562B41DFC09";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F7040370A4C4795EE5606A442810C13C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 772 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"9A1562B41DFC09") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0CD54CE8AB8964293EE42CA28D3D14D0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"9A1562B41DFC09";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0CD54CE8AB8964293EE42CA28D3D14D0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 773 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"9A1562B41DFC09") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"86B9A55141737453F86E20391D87414F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"9A1562B41DFC09";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"86B9A55141737453F86E20391D87414F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 774 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"9A1562B41DFC09") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B763F05941C23BF410FE3FE4CC2CE5C9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"9A1562B41DFC09";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B763F05941C23BF410FE3FE4CC2CE5C9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 775 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"9A1562B41DFC09") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"32BF2F51DDB9E2E21C4AE46FB66942C5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"9A1562B41DFC09";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"32BF2F51DDB9E2E21C4AE46FB66942C5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 776 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"9A1562B41DFC09") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"823E740C76BAA465246CA509BFC20A1B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"9A1562B41DFC09";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"823E740C76BAA465246CA509BFC20A1B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 777 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"9A1562B41DFC09") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3C384CD9456A6665DC11C29B868581F1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"9A1562B41DFC09";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3C384CD9456A6665DC11C29B868581F1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 778 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"9A1562B41DFC09") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0396B8B38E6A384E7AB67172DB27AF4C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"9A1562B41DFC09";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0396B8B38E6A384E7AB67172DB27AF4C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 779 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"9A1562B41DFC09") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9BE1C099AE7A63BC06A867AC00A9DC9C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"9A1562B41DFC09";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9BE1C099AE7A63BC06A867AC00A9DC9C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 780 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"9A1562B41DFC09") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E7D721AC4AC4A8131BDA703B1EDA092B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"9A1562B41DFC09";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E7D721AC4AC4A8131BDA703B1EDA092B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 781 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"9A1562B41DFC09") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E737717752609D172AC132D896A1CF79") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"9A1562B41DFC09";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E737717752609D172AC132D896A1CF79") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 782 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"9A1562B41DFC09") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"34CEE0A1E666C66500838AC8742D07F6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"9A1562B41DFC09";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"34CEE0A1E666C66500838AC8742D07F6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 783 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"9A1562B41DFC09") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F2DBE0BBE6292606A81C3CAA75B13074") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"9A1562B41DFC09";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F2DBE0BBE6292606A81C3CAA75B13074") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 784 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"9A1562B41DFC09") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"74C2B8575B5F101D4BC6130E52AA0EE2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"9A1562B41DFC09";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"74C2B8575B5F101D4BC6130E52AA0EE2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 785 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"9A1562B41DFC09") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DFB96C5053265766FE8A1B017EA6A892") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"9A1562B41DFC09";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DFB96C5053265766FE8A1B017EA6A892") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 786 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"9A1562B41DFC09") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C6DD72A152538CB65A10477B0041C3D2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"9A1562B41DFC09";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C6DD72A152538CB65A10477B0041C3D2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 787 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"9A1562B41DFC09") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"730D88605C87F4706A753E275CC2E4E1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"9A1562B41DFC09";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"730D88605C87F4706A753E275CC2E4E1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 788 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"9A1562B41DFC09") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BD73FFDA80C361AE6CD450EB7FE5D7A3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"9A1562B41DFC09";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BD73FFDA80C361AE6CD450EB7FE5D7A3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 789 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"9A1562B41DFC09") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0788B5EFCA6033080F2D69B32A040CA8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"9A1562B41DFC09";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0788B5EFCA6033080F2D69B32A040CA8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 790 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"9A1562B41DFC09") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A433CEA43311F072DECE4E684A307FAD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"9A1562B41DFC09";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A433CEA43311F072DECE4E684A307FAD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 791 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"9A1562B41DFC09") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FC82BE57DFAE72A7AF447FB03EFA0BC6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"9A1562B41DFC09";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FC82BE57DFAE72A7AF447FB03EFA0BC6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 792 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"9A1562B41DFC09") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C24F0BC455849BC2BFE58BA666F14B49") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"9A1562B41DFC09";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C24F0BC455849BC2BFE58BA666F14B49") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 793 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"9A1562B41DFC09AF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6C940631F6A5A1A8E37CC7155D903810") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"9A1562B41DFC09AF";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6C940631F6A5A1A8E37CC7155D903810") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 794 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"9A1562B41DFC09AF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B27A8634BB75D291DE3C2A6CADB78289") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"9A1562B41DFC09AF";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B27A8634BB75D291DE3C2A6CADB78289") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 795 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"9A1562B41DFC09AF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9352401ADE879E35678BF33C29EFE356") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"9A1562B41DFC09AF";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9352401ADE879E35678BF33C29EFE356") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 796 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"9A1562B41DFC09AF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"37C5B1E06676A3494A398A3FD84E3FC9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"9A1562B41DFC09AF";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"37C5B1E06676A3494A398A3FD84E3FC9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 797 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"9A1562B41DFC09AF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3F4340DF8362F3DB0BBE9A28FB0A42FA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"9A1562B41DFC09AF";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3F4340DF8362F3DB0BBE9A28FB0A42FA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 798 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"9A1562B41DFC09AF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2BD00C53C44701F772A16140137C1850") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"9A1562B41DFC09AF";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2BD00C53C44701F772A16140137C1850") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 799 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"9A1562B41DFC09AF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1FAD1DB0BB9866F3C08964454039F002") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"9A1562B41DFC09AF";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1FAD1DB0BB9866F3C08964454039F002") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 800 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"9A1562B41DFC09AF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"222B6C58A15CC693234FB6B2ACB12D92") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"9A1562B41DFC09AF";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"222B6C58A15CC693234FB6B2ACB12D92") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 801 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"9A1562B41DFC09AF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0FD98DDE5B3EF70326CB51504D40885C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"9A1562B41DFC09AF";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0FD98DDE5B3EF70326CB51504D40885C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 802 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"9A1562B41DFC09AF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3EAA4844A4A1039B827F96C54BE56B1C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"9A1562B41DFC09AF";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3EAA4844A4A1039B827F96C54BE56B1C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 803 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"9A1562B41DFC09AF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CD3629B3B62D87C5223BF99568635413") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"9A1562B41DFC09AF";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CD3629B3B62D87C5223BF99568635413") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 804 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"9A1562B41DFC09AF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F62AC27A99DAF083CE9357EB504306A7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"9A1562B41DFC09AF";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F62AC27A99DAF083CE9357EB504306A7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 805 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"9A1562B41DFC09AF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0DFB8DE29697EDF41517110DF56ED34B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"9A1562B41DFC09AF";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0DFB8DE29697EDF41517110DF56ED34B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 806 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"9A1562B41DFC09AF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8797645B7C6DFD8ED39D1D9665D486D4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"9A1562B41DFC09AF";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8797645B7C6DFD8ED39D1D9665D486D4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 807 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"9A1562B41DFC09AF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B64D31537CDCB2293B0D024BB47F2252") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"9A1562B41DFC09AF";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B64D31537CDCB2293B0D024BB47F2252") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 808 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"9A1562B41DFC09AF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3391EE5BE0A76B3F37B9D9C0CE3A855E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"9A1562B41DFC09AF";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3391EE5BE0A76B3F37B9D9C0CE3A855E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 809 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"9A1562B41DFC09AF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8310B5064BA42DB80F9F98A6C791CD80") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"9A1562B41DFC09AF";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8310B5064BA42DB80F9F98A6C791CD80") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 810 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"9A1562B41DFC09AF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3D168DD37874EFB8F7E2FF34FED6466A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"9A1562B41DFC09AF";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3D168DD37874EFB8F7E2FF34FED6466A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 811 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"9A1562B41DFC09AF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"02B879B9B374B19351454CDDA37468D7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"9A1562B41DFC09AF";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"02B879B9B374B19351454CDDA37468D7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 812 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"9A1562B41DFC09AF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9ACF01939364EA612D5B5A0378FA1B07") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"9A1562B41DFC09AF";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9ACF01939364EA612D5B5A0378FA1B07") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 813 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"9A1562B41DFC09AF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E6F9E0A677DA21CE30294D946689CEB0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"9A1562B41DFC09AF";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E6F9E0A677DA21CE30294D946689CEB0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 814 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"9A1562B41DFC09AF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E619B07D6F7E14CA01320F77EEF208E2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"9A1562B41DFC09AF";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E619B07D6F7E14CA01320F77EEF208E2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 815 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"9A1562B41DFC09AF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"35E021ABDB784FB82B70B7670C7EC06D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"9A1562B41DFC09AF";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"35E021ABDB784FB82B70B7670C7EC06D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 816 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"9A1562B41DFC09AF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F3F521B1DB37AFDB83EF01050DE2F7EF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"9A1562B41DFC09AF";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F3F521B1DB37AFDB83EF01050DE2F7EF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 817 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"9A1562B41DFC09AF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"75EC795D664199C060352EA12AF9C979") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"9A1562B41DFC09AF";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"75EC795D664199C060352EA12AF9C979") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 818 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"9A1562B41DFC09AF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DE97AD5A6E38DEBBD57926AE06F56F09") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"9A1562B41DFC09AF";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DE97AD5A6E38DEBBD57926AE06F56F09") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 819 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"9A1562B41DFC09AF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C7F3B3AB6F4D056B71E37AD478120449") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"9A1562B41DFC09AF";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C7F3B3AB6F4D056B71E37AD478120449") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 820 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"9A1562B41DFC09AF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7223496A61997DAD418603882491237A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"9A1562B41DFC09AF";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7223496A61997DAD418603882491237A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 821 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"9A1562B41DFC09AF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BC5D3ED0BDDDE87347276D4407B61038") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"9A1562B41DFC09AF";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BC5D3ED0BDDDE87347276D4407B61038") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 822 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"9A1562B41DFC09AF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"06A674E5F77EBAD524DE541C5257CB33") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"9A1562B41DFC09AF";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"06A674E5F77EBAD524DE541C5257CB33") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 823 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"9A1562B41DFC09AF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A51D0FAE0E0F79AFF53D73C73263B836") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"9A1562B41DFC09AF";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A51D0FAE0E0F79AFF53D73C73263B836") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 824 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"9A1562B41DFC09AF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FDAC7F5DE2B0FB7A84B7421F46A9CC5D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"9A1562B41DFC09AF";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FDAC7F5DE2B0FB7A84B7421F46A9CC5D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 825 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"9A1562B41DFC09AF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C361CACE689A121F9416B6091EA28CD2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"9A1562B41DFC09AF";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C361CACE689A121F9416B6091EA28CD2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 826 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"9A1562B41DFC09AF6C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E89CD424C0BFB41EE762F0A93B8CA6DA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"9A1562B41DFC09AF6C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E89CD424C0BFB41EE762F0A93B8CA6DA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 827 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"9A1562B41DFC09AF6C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"367254218D6FC727DA221DD0CBAB1C43") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"9A1562B41DFC09AF6C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"367254218D6FC727DA221DD0CBAB1C43") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 828 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"9A1562B41DFC09AF6C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"175A920FE89D8B836395C4804FF37D9C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"9A1562B41DFC09AF6C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"175A920FE89D8B836395C4804FF37D9C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 829 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"9A1562B41DFC09AF6C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B3CD63F5506CB6FF4E27BD83BE52A103") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"9A1562B41DFC09AF6C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B3CD63F5506CB6FF4E27BD83BE52A103") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 830 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"9A1562B41DFC09AF6C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BB4B92CAB578E66D0FA0AD949D16DC30") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"9A1562B41DFC09AF6C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BB4B92CAB578E66D0FA0AD949D16DC30") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 831 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"9A1562B41DFC09AF6C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AFD8DE46F25D144176BF56FC7560869A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"9A1562B41DFC09AF6C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AFD8DE46F25D144176BF56FC7560869A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 832 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"9A1562B41DFC09AF6C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9BA5CFA58D827345C49753F926256EC8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"9A1562B41DFC09AF6C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9BA5CFA58D827345C49753F926256EC8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 833 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"9A1562B41DFC09AF6C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A623BE4D9746D3252751810ECAADB358") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"9A1562B41DFC09AF6C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A623BE4D9746D3252751810ECAADB358") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 834 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"9A1562B41DFC09AF6C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8BD15FCB6D24E2B522D566EC2B5C1696") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"9A1562B41DFC09AF6C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8BD15FCB6D24E2B522D566EC2B5C1696") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 835 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"9A1562B41DFC09AF6C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BAA29A5192BB162D8661A1792DF9F5D6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"9A1562B41DFC09AF6C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BAA29A5192BB162D8661A1792DF9F5D6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 836 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"9A1562B41DFC09AF6C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"493EFBA6803792732625CE290E7FCAD9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"9A1562B41DFC09AF6C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"493EFBA6803792732625CE290E7FCAD9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 837 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"9A1562B41DFC09AF6C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7222106FAFC0E535CA8D6057365F986D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"9A1562B41DFC09AF6C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7222106FAFC0E535CA8D6057365F986D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 838 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"9A1562B41DFC09AF6C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"89F35FF7A08DF842110926B193724D81") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"9A1562B41DFC09AF6C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"89F35FF7A08DF842110926B193724D81") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 839 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"9A1562B41DFC09AF6C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"039FB64E4A77E838D7832A2A03C8181E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"9A1562B41DFC09AF6C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"039FB64E4A77E838D7832A2A03C8181E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 840 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"9A1562B41DFC09AF6C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3245E3464AC6A79F3F1335F7D263BC98") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"9A1562B41DFC09AF6C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3245E3464AC6A79F3F1335F7D263BC98") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 841 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"9A1562B41DFC09AF6C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B7993C4ED6BD7E8933A7EE7CA8261B94") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"9A1562B41DFC09AF6C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B7993C4ED6BD7E8933A7EE7CA8261B94") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 842 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"9A1562B41DFC09AF6C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"071867137DBE380E0B81AF1AA18D534A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"9A1562B41DFC09AF6C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"071867137DBE380E0B81AF1AA18D534A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 843 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"9A1562B41DFC09AF6C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B91E5FC64E6EFA0EF3FCC88898CAD8A0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"9A1562B41DFC09AF6C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B91E5FC64E6EFA0EF3FCC88898CAD8A0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 844 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"9A1562B41DFC09AF6C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"86B0ABAC856EA425555B7B61C568F61D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"9A1562B41DFC09AF6C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"86B0ABAC856EA425555B7B61C568F61D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 845 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"9A1562B41DFC09AF6C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1EC7D386A57EFFD729456DBF1EE685CD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"9A1562B41DFC09AF6C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1EC7D386A57EFFD729456DBF1EE685CD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 846 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"9A1562B41DFC09AF6C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"62F132B341C0347834377A280095507A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"9A1562B41DFC09AF6C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"62F132B341C0347834377A280095507A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 847 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"9A1562B41DFC09AF6C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"621162685964017C052C38CB88EE9628") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"9A1562B41DFC09AF6C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"621162685964017C052C38CB88EE9628") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 848 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"9A1562B41DFC09AF6C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B1E8F3BEED625A0E2F6E80DB6A625EA7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"9A1562B41DFC09AF6C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B1E8F3BEED625A0E2F6E80DB6A625EA7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 849 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"9A1562B41DFC09AF6C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"77FDF3A4ED2DBA6D87F136B96BFE6925") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"9A1562B41DFC09AF6C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"77FDF3A4ED2DBA6D87F136B96BFE6925") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 850 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"9A1562B41DFC09AF6C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F1E4AB48505B8C76642B191D4CE557B3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"9A1562B41DFC09AF6C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F1E4AB48505B8C76642B191D4CE557B3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 851 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"9A1562B41DFC09AF6C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5A9F7F4F5822CB0DD167111260E9F1C3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"9A1562B41DFC09AF6C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5A9F7F4F5822CB0DD167111260E9F1C3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 852 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"9A1562B41DFC09AF6C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"43FB61BE595710DD75FD4D681E0E9A83") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"9A1562B41DFC09AF6C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"43FB61BE595710DD75FD4D681E0E9A83") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 853 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"9A1562B41DFC09AF6C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F62B9B7F5783681B45983434428DBDB0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"9A1562B41DFC09AF6C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F62B9B7F5783681B45983434428DBDB0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 854 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"9A1562B41DFC09AF6C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3855ECC58BC7FDC543395AF861AA8EF2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"9A1562B41DFC09AF6C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3855ECC58BC7FDC543395AF861AA8EF2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 855 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"9A1562B41DFC09AF6C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"82AEA6F0C164AF6320C063A0344B55F9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"9A1562B41DFC09AF6C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"82AEA6F0C164AF6320C063A0344B55F9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 856 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"9A1562B41DFC09AF6C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2115DDBB38156C19F123447B547F26FC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"9A1562B41DFC09AF6C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2115DDBB38156C19F123447B547F26FC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 857 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"9A1562B41DFC09AF6C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"79A4AD48D4AAEECC80A975A320B55297") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"9A1562B41DFC09AF6C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"79A4AD48D4AAEECC80A975A320B55297") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 858 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"9A1562B41DFC09AF6C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"476918DB5E8007A9900881B578BE1218") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"9A1562B41DFC09AF6C";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"476918DB5E8007A9900881B578BE1218") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 859 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"9A1562B41DFC09AF6C55") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8E0A7DCC7DB2278F218335D89FFDE741") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"9A1562B41DFC09AF6C55";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8E0A7DCC7DB2278F218335D89FFDE741") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 860 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"9A1562B41DFC09AF6C55") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"50E4FDC9306254B61CC3D8A16FDA5DD8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"9A1562B41DFC09AF6C55";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"50E4FDC9306254B61CC3D8A16FDA5DD8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 861 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"9A1562B41DFC09AF6C55") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"71CC3BE755901812A57401F1EB823C07") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"9A1562B41DFC09AF6C55";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"71CC3BE755901812A57401F1EB823C07") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 862 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"9A1562B41DFC09AF6C55") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D55BCA1DED61256E88C678F21A23E098") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"9A1562B41DFC09AF6C55";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D55BCA1DED61256E88C678F21A23E098") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 863 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"9A1562B41DFC09AF6C55") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DDDD3B22087575FCC94168E539679DAB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"9A1562B41DFC09AF6C55";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DDDD3B22087575FCC94168E539679DAB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 864 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"9A1562B41DFC09AF6C55") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C94E77AE4F5087D0B05E938DD111C701") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"9A1562B41DFC09AF6C55";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C94E77AE4F5087D0B05E938DD111C701") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 865 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"9A1562B41DFC09AF6C55") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FD33664D308FE0D40276968882542F53") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"9A1562B41DFC09AF6C55";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FD33664D308FE0D40276968882542F53") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 866 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"9A1562B41DFC09AF6C55") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C0B517A52A4B40B4E1B0447F6EDCF2C3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"9A1562B41DFC09AF6C55";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C0B517A52A4B40B4E1B0447F6EDCF2C3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 867 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"9A1562B41DFC09AF6C55") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"ED47F623D0297124E434A39D8F2D570D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"9A1562B41DFC09AF6C55";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"ED47F623D0297124E434A39D8F2D570D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 868 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"9A1562B41DFC09AF6C55") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DC3433B92FB685BC408064088988B44D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"9A1562B41DFC09AF6C55";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DC3433B92FB685BC408064088988B44D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 869 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"9A1562B41DFC09AF6C55") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2FA8524E3D3A01E2E0C40B58AA0E8B42") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"9A1562B41DFC09AF6C55";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2FA8524E3D3A01E2E0C40B58AA0E8B42") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 870 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"9A1562B41DFC09AF6C55") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"14B4B98712CD76A40C6CA526922ED9F6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"9A1562B41DFC09AF6C55";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"14B4B98712CD76A40C6CA526922ED9F6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 871 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"9A1562B41DFC09AF6C55") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EF65F61F1D806BD3D7E8E3C037030C1A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"9A1562B41DFC09AF6C55";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EF65F61F1D806BD3D7E8E3C037030C1A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 872 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"9A1562B41DFC09AF6C55") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"65091FA6F77A7BA91162EF5BA7B95985") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"9A1562B41DFC09AF6C55";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"65091FA6F77A7BA91162EF5BA7B95985") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 873 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"9A1562B41DFC09AF6C55") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"54D34AAEF7CB340EF9F2F0867612FD03") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"9A1562B41DFC09AF6C55";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"54D34AAEF7CB340EF9F2F0867612FD03") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 874 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"9A1562B41DFC09AF6C55") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D10F95A66BB0ED18F5462B0D0C575A0F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"9A1562B41DFC09AF6C55";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D10F95A66BB0ED18F5462B0D0C575A0F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 875 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"9A1562B41DFC09AF6C55") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"618ECEFBC0B3AB9FCD606A6B05FC12D1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"9A1562B41DFC09AF6C55";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"618ECEFBC0B3AB9FCD606A6B05FC12D1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 876 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"9A1562B41DFC09AF6C55") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DF88F62EF363699F351D0DF93CBB993B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"9A1562B41DFC09AF6C55";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DF88F62EF363699F351D0DF93CBB993B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 877 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"9A1562B41DFC09AF6C55") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E0260244386337B493BABE106119B786") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"9A1562B41DFC09AF6C55";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E0260244386337B493BABE106119B786") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 878 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"9A1562B41DFC09AF6C55") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"78517A6E18736C46EFA4A8CEBA97C456") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"9A1562B41DFC09AF6C55";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"78517A6E18736C46EFA4A8CEBA97C456") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 879 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"9A1562B41DFC09AF6C55") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"04679B5BFCCDA7E9F2D6BF59A4E411E1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"9A1562B41DFC09AF6C55";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"04679B5BFCCDA7E9F2D6BF59A4E411E1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 880 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"9A1562B41DFC09AF6C55") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0487CB80E46992EDC3CDFDBA2C9FD7B3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"9A1562B41DFC09AF6C55";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0487CB80E46992EDC3CDFDBA2C9FD7B3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 881 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"9A1562B41DFC09AF6C55") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D77E5A56506FC99FE98F45AACE131F3C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"9A1562B41DFC09AF6C55";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D77E5A56506FC99FE98F45AACE131F3C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 882 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"9A1562B41DFC09AF6C55") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"116B5A4C502029FC4110F3C8CF8F28BE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"9A1562B41DFC09AF6C55";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"116B5A4C502029FC4110F3C8CF8F28BE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 883 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"9A1562B41DFC09AF6C55") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"977202A0ED561FE7A2CADC6CE8941628") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"9A1562B41DFC09AF6C55";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"977202A0ED561FE7A2CADC6CE8941628") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 884 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"9A1562B41DFC09AF6C55") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3C09D6A7E52F589C1786D463C498B058") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"9A1562B41DFC09AF6C55";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3C09D6A7E52F589C1786D463C498B058") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 885 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"9A1562B41DFC09AF6C55") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"256DC856E45A834CB31C8819BA7FDB18") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"9A1562B41DFC09AF6C55";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"256DC856E45A834CB31C8819BA7FDB18") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 886 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"9A1562B41DFC09AF6C55") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"90BD3297EA8EFB8A8379F145E6FCFC2B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"9A1562B41DFC09AF6C55";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"90BD3297EA8EFB8A8379F145E6FCFC2B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 887 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"9A1562B41DFC09AF6C55") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5EC3452D36CA6E5485D89F89C5DBCF69") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"9A1562B41DFC09AF6C55";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5EC3452D36CA6E5485D89F89C5DBCF69") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 888 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"9A1562B41DFC09AF6C55") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E4380F187C693CF2E621A6D1903A1462") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"9A1562B41DFC09AF6C55";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E4380F187C693CF2E621A6D1903A1462") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 889 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"9A1562B41DFC09AF6C55") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"478374538518FF8837C2810AF00E6767") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"9A1562B41DFC09AF6C55";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"478374538518FF8837C2810AF00E6767") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 890 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"9A1562B41DFC09AF6C55") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1F3204A069A77D5D4648B0D284C4130C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"9A1562B41DFC09AF6C55";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1F3204A069A77D5D4648B0D284C4130C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 891 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"9A1562B41DFC09AF6C55") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"21FFB133E38D943856E944C4DCCF5383") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"9A1562B41DFC09AF6C55";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"21FFB133E38D943856E944C4DCCF5383") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 892 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"9A1562B41DFC09AF6C55EC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BA5AC4191A6ACBC8BAD461960E1FBB9A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"9A1562B41DFC09AF6C55EC";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BA5AC4191A6ACBC8BAD461960E1FBB9A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 893 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"9A1562B41DFC09AF6C55EC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"64B4441C57BAB8F187948CEFFE380103") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"9A1562B41DFC09AF6C55EC";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"64B4441C57BAB8F187948CEFFE380103") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 894 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"9A1562B41DFC09AF6C55EC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"459C82323248F4553E2355BF7A6060DC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"9A1562B41DFC09AF6C55EC";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"459C82323248F4553E2355BF7A6060DC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 895 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"9A1562B41DFC09AF6C55EC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E10B73C88AB9C92913912CBC8BC1BC43") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"9A1562B41DFC09AF6C55EC";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E10B73C88AB9C92913912CBC8BC1BC43") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 896 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"9A1562B41DFC09AF6C55EC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E98D82F76FAD99BB52163CABA885C170") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"9A1562B41DFC09AF6C55EC";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E98D82F76FAD99BB52163CABA885C170") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 897 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"9A1562B41DFC09AF6C55EC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FD1ECE7B28886B972B09C7C340F39BDA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"9A1562B41DFC09AF6C55EC";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FD1ECE7B28886B972B09C7C340F39BDA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 898 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"9A1562B41DFC09AF6C55EC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C963DF9857570C939921C2C613B67388") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"9A1562B41DFC09AF6C55EC";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C963DF9857570C939921C2C613B67388") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 899 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"9A1562B41DFC09AF6C55EC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F4E5AE704D93ACF37AE71031FF3EAE18") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"9A1562B41DFC09AF6C55EC";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F4E5AE704D93ACF37AE71031FF3EAE18") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 900 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"9A1562B41DFC09AF6C55EC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D9174FF6B7F19D637F63F7D31ECF0BD6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"9A1562B41DFC09AF6C55EC";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D9174FF6B7F19D637F63F7D31ECF0BD6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 901 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"9A1562B41DFC09AF6C55EC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E8648A6C486E69FBDBD73046186AE896") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"9A1562B41DFC09AF6C55EC";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E8648A6C486E69FBDBD73046186AE896") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 902 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"9A1562B41DFC09AF6C55EC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1BF8EB9B5AE2EDA57B935F163BECD799") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"9A1562B41DFC09AF6C55EC";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1BF8EB9B5AE2EDA57B935F163BECD799") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 903 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"9A1562B41DFC09AF6C55EC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"20E4005275159AE3973BF16803CC852D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"9A1562B41DFC09AF6C55EC";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"20E4005275159AE3973BF16803CC852D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 904 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"9A1562B41DFC09AF6C55EC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DB354FCA7A5887944CBFB78EA6E150C1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"9A1562B41DFC09AF6C55EC";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DB354FCA7A5887944CBFB78EA6E150C1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 905 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"9A1562B41DFC09AF6C55EC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5159A67390A297EE8A35BB15365B055E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"9A1562B41DFC09AF6C55EC";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5159A67390A297EE8A35BB15365B055E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 906 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"9A1562B41DFC09AF6C55EC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6083F37B9013D84962A5A4C8E7F0A1D8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"9A1562B41DFC09AF6C55EC";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6083F37B9013D84962A5A4C8E7F0A1D8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 907 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"9A1562B41DFC09AF6C55EC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E55F2C730C68015F6E117F439DB506D4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"9A1562B41DFC09AF6C55EC";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E55F2C730C68015F6E117F439DB506D4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 908 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"9A1562B41DFC09AF6C55EC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"55DE772EA76B47D856373E25941E4E0A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"9A1562B41DFC09AF6C55EC";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"55DE772EA76B47D856373E25941E4E0A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 909 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"9A1562B41DFC09AF6C55EC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EBD84FFB94BB85D8AE4A59B7AD59C5E0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"9A1562B41DFC09AF6C55EC";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EBD84FFB94BB85D8AE4A59B7AD59C5E0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 910 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"9A1562B41DFC09AF6C55EC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D476BB915FBBDBF308EDEA5EF0FBEB5D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"9A1562B41DFC09AF6C55EC";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D476BB915FBBDBF308EDEA5EF0FBEB5D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 911 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"9A1562B41DFC09AF6C55EC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4C01C3BB7FAB800174F3FC802B75988D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"9A1562B41DFC09AF6C55EC";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4C01C3BB7FAB800174F3FC802B75988D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 912 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"9A1562B41DFC09AF6C55EC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3037228E9B154BAE6981EB1735064D3A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"9A1562B41DFC09AF6C55EC";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3037228E9B154BAE6981EB1735064D3A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 913 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"9A1562B41DFC09AF6C55EC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"30D7725583B17EAA589AA9F4BD7D8B68") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"9A1562B41DFC09AF6C55EC";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"30D7725583B17EAA589AA9F4BD7D8B68") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 914 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"9A1562B41DFC09AF6C55EC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E32EE38337B725D872D811E45FF143E7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"9A1562B41DFC09AF6C55EC";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E32EE38337B725D872D811E45FF143E7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 915 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"9A1562B41DFC09AF6C55EC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"253BE39937F8C5BBDA47A7865E6D7465") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"9A1562B41DFC09AF6C55EC";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"253BE39937F8C5BBDA47A7865E6D7465") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 916 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"9A1562B41DFC09AF6C55EC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A322BB758A8EF3A0399D882279764AF3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"9A1562B41DFC09AF6C55EC";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A322BB758A8EF3A0399D882279764AF3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 917 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"9A1562B41DFC09AF6C55EC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"08596F7282F7B4DB8CD1802D557AEC83") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"9A1562B41DFC09AF6C55EC";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"08596F7282F7B4DB8CD1802D557AEC83") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 918 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"9A1562B41DFC09AF6C55EC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"113D718383826F0B284BDC572B9D87C3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"9A1562B41DFC09AF6C55EC";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"113D718383826F0B284BDC572B9D87C3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 919 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"9A1562B41DFC09AF6C55EC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A4ED8B428D5617CD182EA50B771EA0F0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"9A1562B41DFC09AF6C55EC";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A4ED8B428D5617CD182EA50B771EA0F0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 920 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"9A1562B41DFC09AF6C55EC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6A93FCF8511282131E8FCBC7543993B2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"9A1562B41DFC09AF6C55EC";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6A93FCF8511282131E8FCBC7543993B2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 921 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"9A1562B41DFC09AF6C55EC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D068B6CD1BB1D0B57D76F29F01D848B9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"9A1562B41DFC09AF6C55EC";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D068B6CD1BB1D0B57D76F29F01D848B9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 922 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"9A1562B41DFC09AF6C55EC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"73D3CD86E2C013CFAC95D54461EC3BBC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"9A1562B41DFC09AF6C55EC";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"73D3CD86E2C013CFAC95D54461EC3BBC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 923 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"9A1562B41DFC09AF6C55EC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2B62BD750E7F911ADD1FE49C15264FD7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"9A1562B41DFC09AF6C55EC";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2B62BD750E7F911ADD1FE49C15264FD7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 924 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"9A1562B41DFC09AF6C55EC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"15AF08E68455787FCDBE108A4D2D0F58") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"9A1562B41DFC09AF6C55EC";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"15AF08E68455787FCDBE108A4D2D0F58") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 925 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"9A1562B41DFC09AF6C55ECD1") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4247C5A2F9FDF576BB4BF69269B9DCA3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"9A1562B41DFC09AF6C55ECD1";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4247C5A2F9FDF576BB4BF69269B9DCA3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 926 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"9A1562B41DFC09AF6C55ECD1") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9CA945A7B42D864F860B1BEB999E663A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"9A1562B41DFC09AF6C55ECD1";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9CA945A7B42D864F860B1BEB999E663A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 927 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"9A1562B41DFC09AF6C55ECD1") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BD818389D1DFCAEB3FBCC2BB1DC607E5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"9A1562B41DFC09AF6C55ECD1";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BD818389D1DFCAEB3FBCC2BB1DC607E5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 928 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"9A1562B41DFC09AF6C55ECD1") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"19167273692EF797120EBBB8EC67DB7A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"9A1562B41DFC09AF6C55ECD1";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"19167273692EF797120EBBB8EC67DB7A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 929 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"9A1562B41DFC09AF6C55ECD1") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1190834C8C3AA7055389ABAFCF23A649") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"9A1562B41DFC09AF6C55ECD1";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1190834C8C3AA7055389ABAFCF23A649") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 930 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"9A1562B41DFC09AF6C55ECD1") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0503CFC0CB1F55292A9650C72755FCE3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"9A1562B41DFC09AF6C55ECD1";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0503CFC0CB1F55292A9650C72755FCE3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 931 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"9A1562B41DFC09AF6C55ECD1") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"317EDE23B4C0322D98BE55C2741014B1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"9A1562B41DFC09AF6C55ECD1";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"317EDE23B4C0322D98BE55C2741014B1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 932 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"9A1562B41DFC09AF6C55ECD1") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0CF8AFCBAE04924D7B7887359898C921") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"9A1562B41DFC09AF6C55ECD1";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0CF8AFCBAE04924D7B7887359898C921") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 933 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"9A1562B41DFC09AF6C55ECD1") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"210A4E4D5466A3DD7EFC60D779696CEF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"9A1562B41DFC09AF6C55ECD1";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"210A4E4D5466A3DD7EFC60D779696CEF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 934 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"9A1562B41DFC09AF6C55ECD1") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"10798BD7ABF95745DA48A7427FCC8FAF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"9A1562B41DFC09AF6C55ECD1";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"10798BD7ABF95745DA48A7427FCC8FAF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 935 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"9A1562B41DFC09AF6C55ECD1") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E3E5EA20B975D31B7A0CC8125C4AB0A0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"9A1562B41DFC09AF6C55ECD1";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E3E5EA20B975D31B7A0CC8125C4AB0A0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 936 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"9A1562B41DFC09AF6C55ECD1") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D8F901E99682A45D96A4666C646AE214") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"9A1562B41DFC09AF6C55ECD1";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D8F901E99682A45D96A4666C646AE214") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 937 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"9A1562B41DFC09AF6C55ECD1") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"23284E7199CFB92A4D20208AC14737F8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"9A1562B41DFC09AF6C55ECD1";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"23284E7199CFB92A4D20208AC14737F8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 938 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"9A1562B41DFC09AF6C55ECD1") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A944A7C87335A9508BAA2C1151FD6267") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"9A1562B41DFC09AF6C55ECD1";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A944A7C87335A9508BAA2C1151FD6267") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 939 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"9A1562B41DFC09AF6C55ECD1") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"989EF2C07384E6F7633A33CC8056C6E1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"9A1562B41DFC09AF6C55ECD1";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"989EF2C07384E6F7633A33CC8056C6E1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 940 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"9A1562B41DFC09AF6C55ECD1") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1D422DC8EFFF3FE16F8EE847FA1361ED") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"9A1562B41DFC09AF6C55ECD1";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1D422DC8EFFF3FE16F8EE847FA1361ED") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 941 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"9A1562B41DFC09AF6C55ECD1") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"ADC3769544FC796657A8A921F3B82933") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"9A1562B41DFC09AF6C55ECD1";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"ADC3769544FC796657A8A921F3B82933") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 942 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"9A1562B41DFC09AF6C55ECD1") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"13C54E40772CBB66AFD5CEB3CAFFA2D9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"9A1562B41DFC09AF6C55ECD1";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"13C54E40772CBB66AFD5CEB3CAFFA2D9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 943 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"9A1562B41DFC09AF6C55ECD1") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2C6BBA2ABC2CE54D09727D5A975D8C64") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"9A1562B41DFC09AF6C55ECD1";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2C6BBA2ABC2CE54D09727D5A975D8C64") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 944 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"9A1562B41DFC09AF6C55ECD1") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B41CC2009C3CBEBF756C6B844CD3FFB4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"9A1562B41DFC09AF6C55ECD1";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B41CC2009C3CBEBF756C6B844CD3FFB4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 945 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"9A1562B41DFC09AF6C55ECD1") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C82A233578827510681E7C1352A02A03") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"9A1562B41DFC09AF6C55ECD1";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C82A233578827510681E7C1352A02A03") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 946 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"9A1562B41DFC09AF6C55ECD1") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C8CA73EE6026401459053EF0DADBEC51") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"9A1562B41DFC09AF6C55ECD1";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C8CA73EE6026401459053EF0DADBEC51") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 947 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"9A1562B41DFC09AF6C55ECD1") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1B33E238D4201B66734786E0385724DE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"9A1562B41DFC09AF6C55ECD1";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1B33E238D4201B66734786E0385724DE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 948 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"9A1562B41DFC09AF6C55ECD1") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DD26E222D46FFB05DBD8308239CB135C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"9A1562B41DFC09AF6C55ECD1";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DD26E222D46FFB05DBD8308239CB135C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 949 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"9A1562B41DFC09AF6C55ECD1") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5B3FBACE6919CD1E38021F261ED02DCA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"9A1562B41DFC09AF6C55ECD1";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5B3FBACE6919CD1E38021F261ED02DCA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 950 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"9A1562B41DFC09AF6C55ECD1") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F0446EC961608A658D4E172932DC8BBA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"9A1562B41DFC09AF6C55ECD1";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F0446EC961608A658D4E172932DC8BBA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 951 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"9A1562B41DFC09AF6C55ECD1") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E9207038601551B529D44B534C3BE0FA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"9A1562B41DFC09AF6C55ECD1";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E9207038601551B529D44B534C3BE0FA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 952 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"9A1562B41DFC09AF6C55ECD1") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5CF08AF96EC1297319B1320F10B8C7C9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"9A1562B41DFC09AF6C55ECD1";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5CF08AF96EC1297319B1320F10B8C7C9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 953 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"9A1562B41DFC09AF6C55ECD1") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"928EFD43B285BCAD1F105CC3339FF48B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"9A1562B41DFC09AF6C55ECD1";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"928EFD43B285BCAD1F105CC3339FF48B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 954 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"9A1562B41DFC09AF6C55ECD1") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2875B776F826EE0B7CE9659B667E2F80") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"9A1562B41DFC09AF6C55ECD1";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2875B776F826EE0B7CE9659B667E2F80") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 955 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"9A1562B41DFC09AF6C55ECD1") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8BCECC3D01572D71AD0A4240064A5C85") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"9A1562B41DFC09AF6C55ECD1";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8BCECC3D01572D71AD0A4240064A5C85") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 956 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"9A1562B41DFC09AF6C55ECD1") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D37FBCCEEDE8AFA4DC807398728028EE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"9A1562B41DFC09AF6C55ECD1";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D37FBCCEEDE8AFA4DC807398728028EE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 957 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"9A1562B41DFC09AF6C55ECD1") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EDB2095D67C246C1CC21878E2A8B6861") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"9A1562B41DFC09AF6C55ECD1";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EDB2095D67C246C1CC21878E2A8B6861") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 958 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"9A1562B41DFC09AF6C55ECD14D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"152914CF4E5B47E598246EED8D33CF87") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"9A1562B41DFC09AF6C55ECD14D";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"152914CF4E5B47E598246EED8D33CF87") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 959 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"9A1562B41DFC09AF6C55ECD14D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CBC794CA038B34DCA56483947D14751E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"9A1562B41DFC09AF6C55ECD14D";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CBC794CA038B34DCA56483947D14751E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 960 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"9A1562B41DFC09AF6C55ECD14D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EAEF52E4667978781CD35AC4F94C14C1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"9A1562B41DFC09AF6C55ECD14D";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EAEF52E4667978781CD35AC4F94C14C1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 961 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"9A1562B41DFC09AF6C55ECD14D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4E78A31EDE884504316123C708EDC85E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"9A1562B41DFC09AF6C55ECD14D";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4E78A31EDE884504316123C708EDC85E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 962 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"9A1562B41DFC09AF6C55ECD14D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"46FE52213B9C159670E633D02BA9B56D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"9A1562B41DFC09AF6C55ECD14D";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"46FE52213B9C159670E633D02BA9B56D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 963 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"9A1562B41DFC09AF6C55ECD14D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"526D1EAD7CB9E7BA09F9C8B8C3DFEFC7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"9A1562B41DFC09AF6C55ECD14D";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"526D1EAD7CB9E7BA09F9C8B8C3DFEFC7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 964 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"9A1562B41DFC09AF6C55ECD14D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"66100F4E036680BEBBD1CDBD909A0795") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"9A1562B41DFC09AF6C55ECD14D";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"66100F4E036680BEBBD1CDBD909A0795") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 965 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"9A1562B41DFC09AF6C55ECD14D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5B967EA619A220DE58171F4A7C12DA05") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"9A1562B41DFC09AF6C55ECD14D";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5B967EA619A220DE58171F4A7C12DA05") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 966 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"9A1562B41DFC09AF6C55ECD14D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"76649F20E3C0114E5D93F8A89DE37FCB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"9A1562B41DFC09AF6C55ECD14D";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"76649F20E3C0114E5D93F8A89DE37FCB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 967 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"9A1562B41DFC09AF6C55ECD14D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"47175ABA1C5FE5D6F9273F3D9B469C8B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"9A1562B41DFC09AF6C55ECD14D";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"47175ABA1C5FE5D6F9273F3D9B469C8B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 968 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"9A1562B41DFC09AF6C55ECD14D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B48B3B4D0ED361885963506DB8C0A384") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"9A1562B41DFC09AF6C55ECD14D";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B48B3B4D0ED361885963506DB8C0A384") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 969 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"9A1562B41DFC09AF6C55ECD14D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8F97D084212416CEB5CBFE1380E0F130") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"9A1562B41DFC09AF6C55ECD14D";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8F97D084212416CEB5CBFE1380E0F130") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 970 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"9A1562B41DFC09AF6C55ECD14D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"74469F1C2E690BB96E4FB8F525CD24DC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"9A1562B41DFC09AF6C55ECD14D";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"74469F1C2E690BB96E4FB8F525CD24DC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 971 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"9A1562B41DFC09AF6C55ECD14D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FE2A76A5C4931BC3A8C5B46EB5777143") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"9A1562B41DFC09AF6C55ECD14D";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FE2A76A5C4931BC3A8C5B46EB5777143") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 972 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"9A1562B41DFC09AF6C55ECD14D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CFF023ADC42254644055ABB364DCD5C5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"9A1562B41DFC09AF6C55ECD14D";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CFF023ADC42254644055ABB364DCD5C5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 973 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"9A1562B41DFC09AF6C55ECD14D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4A2CFCA558598D724CE170381E9972C9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"9A1562B41DFC09AF6C55ECD14D";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4A2CFCA558598D724CE170381E9972C9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 974 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"9A1562B41DFC09AF6C55ECD14D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FAADA7F8F35ACBF574C7315E17323A17") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"9A1562B41DFC09AF6C55ECD14D";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FAADA7F8F35ACBF574C7315E17323A17") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 975 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"9A1562B41DFC09AF6C55ECD14D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"44AB9F2DC08A09F58CBA56CC2E75B1FD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"9A1562B41DFC09AF6C55ECD14D";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"44AB9F2DC08A09F58CBA56CC2E75B1FD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 976 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"9A1562B41DFC09AF6C55ECD14D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7B056B470B8A57DE2A1DE52573D79F40") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"9A1562B41DFC09AF6C55ECD14D";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7B056B470B8A57DE2A1DE52573D79F40") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 977 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"9A1562B41DFC09AF6C55ECD14D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E372136D2B9A0C2C5603F3FBA859EC90") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"9A1562B41DFC09AF6C55ECD14D";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E372136D2B9A0C2C5603F3FBA859EC90") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 978 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"9A1562B41DFC09AF6C55ECD14D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9F44F258CF24C7834B71E46CB62A3927") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"9A1562B41DFC09AF6C55ECD14D";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9F44F258CF24C7834B71E46CB62A3927") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 979 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"9A1562B41DFC09AF6C55ECD14D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9FA4A283D780F2877A6AA68F3E51FF75") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"9A1562B41DFC09AF6C55ECD14D";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9FA4A283D780F2877A6AA68F3E51FF75") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 980 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"9A1562B41DFC09AF6C55ECD14D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4C5D33556386A9F550281E9FDCDD37FA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"9A1562B41DFC09AF6C55ECD14D";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4C5D33556386A9F550281E9FDCDD37FA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 981 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"9A1562B41DFC09AF6C55ECD14D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8A48334F63C94996F8B7A8FDDD410078") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"9A1562B41DFC09AF6C55ECD14D";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8A48334F63C94996F8B7A8FDDD410078") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 982 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"9A1562B41DFC09AF6C55ECD14D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0C516BA3DEBF7F8D1B6D8759FA5A3EEE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"9A1562B41DFC09AF6C55ECD14D";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0C516BA3DEBF7F8D1B6D8759FA5A3EEE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 983 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"9A1562B41DFC09AF6C55ECD14D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A72ABFA4D6C638F6AE218F56D656989E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"9A1562B41DFC09AF6C55ECD14D";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A72ABFA4D6C638F6AE218F56D656989E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 984 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"9A1562B41DFC09AF6C55ECD14D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BE4EA155D7B3E3260ABBD32CA8B1F3DE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"9A1562B41DFC09AF6C55ECD14D";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BE4EA155D7B3E3260ABBD32CA8B1F3DE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 985 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"9A1562B41DFC09AF6C55ECD14D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0B9E5B94D9679BE03ADEAA70F432D4ED") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"9A1562B41DFC09AF6C55ECD14D";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0B9E5B94D9679BE03ADEAA70F432D4ED") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 986 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"9A1562B41DFC09AF6C55ECD14D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C5E02C2E05230E3E3C7FC4BCD715E7AF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"9A1562B41DFC09AF6C55ECD14D";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C5E02C2E05230E3E3C7FC4BCD715E7AF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 987 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"9A1562B41DFC09AF6C55ECD14D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7F1B661B4F805C985F86FDE482F43CA4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"9A1562B41DFC09AF6C55ECD14D";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7F1B661B4F805C985F86FDE482F43CA4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 988 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"9A1562B41DFC09AF6C55ECD14D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DCA01D50B6F19FE28E65DA3FE2C04FA1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"9A1562B41DFC09AF6C55ECD14D";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DCA01D50B6F19FE28E65DA3FE2C04FA1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 989 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"9A1562B41DFC09AF6C55ECD14D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"84116DA35A4E1D37FFEFEBE7960A3BCA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"9A1562B41DFC09AF6C55ECD14D";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"84116DA35A4E1D37FFEFEBE7960A3BCA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 990 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"9A1562B41DFC09AF6C55ECD14D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BADCD830D064F452EF4E1FF1CE017B45") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"9A1562B41DFC09AF6C55ECD14D";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BADCD830D064F452EF4E1FF1CE017B45") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 991 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"9A1562B41DFC09AF6C55ECD14D3E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"270B7FF2607452FEBD7E7743B3A32D84") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"9A1562B41DFC09AF6C55ECD14D3E";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"270B7FF2607452FEBD7E7743B3A32D84") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 992 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"9A1562B41DFC09AF6C55ECD14D3E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F9E5FFF72DA421C7803E9A3A4384971D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"9A1562B41DFC09AF6C55ECD14D3E";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F9E5FFF72DA421C7803E9A3A4384971D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 993 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"9A1562B41DFC09AF6C55ECD14D3E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D8CD39D948566D633989436AC7DCF6C2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"9A1562B41DFC09AF6C55ECD14D3E";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D8CD39D948566D633989436AC7DCF6C2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 994 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"9A1562B41DFC09AF6C55ECD14D3E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7C5AC823F0A7501F143B3A69367D2A5D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"9A1562B41DFC09AF6C55ECD14D3E";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7C5AC823F0A7501F143B3A69367D2A5D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 995 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"9A1562B41DFC09AF6C55ECD14D3E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"74DC391C15B3008D55BC2A7E1539576E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"9A1562B41DFC09AF6C55ECD14D3E";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"74DC391C15B3008D55BC2A7E1539576E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 996 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"9A1562B41DFC09AF6C55ECD14D3E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"604F75905296F2A12CA3D116FD4F0DC4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"9A1562B41DFC09AF6C55ECD14D3E";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"604F75905296F2A12CA3D116FD4F0DC4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 997 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"9A1562B41DFC09AF6C55ECD14D3E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"543264732D4995A59E8BD413AE0AE596") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"9A1562B41DFC09AF6C55ECD14D3E";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"543264732D4995A59E8BD413AE0AE596") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 998 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"9A1562B41DFC09AF6C55ECD14D3E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"69B4159B378D35C57D4D06E442823806") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"9A1562B41DFC09AF6C55ECD14D3E";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"69B4159B378D35C57D4D06E442823806") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 999 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"9A1562B41DFC09AF6C55ECD14D3E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4446F41DCDEF045578C9E106A3739DC8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"9A1562B41DFC09AF6C55ECD14D3E";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4446F41DCDEF045578C9E106A3739DC8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1000 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"9A1562B41DFC09AF6C55ECD14D3E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"753531873270F0CDDC7D2693A5D67E88") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"9A1562B41DFC09AF6C55ECD14D3E";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"753531873270F0CDDC7D2693A5D67E88") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1001 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"9A1562B41DFC09AF6C55ECD14D3E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"86A9507020FC74937C3949C386504187") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"9A1562B41DFC09AF6C55ECD14D3E";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"86A9507020FC74937C3949C386504187") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1002 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"9A1562B41DFC09AF6C55ECD14D3E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BDB5BBB90F0B03D59091E7BDBE701333") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"9A1562B41DFC09AF6C55ECD14D3E";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BDB5BBB90F0B03D59091E7BDBE701333") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1003 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"9A1562B41DFC09AF6C55ECD14D3E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4664F42100461EA24B15A15B1B5DC6DF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"9A1562B41DFC09AF6C55ECD14D3E";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4664F42100461EA24B15A15B1B5DC6DF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1004 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"9A1562B41DFC09AF6C55ECD14D3E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CC081D98EABC0ED88D9FADC08BE79340") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"9A1562B41DFC09AF6C55ECD14D3E";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CC081D98EABC0ED88D9FADC08BE79340") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1005 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"9A1562B41DFC09AF6C55ECD14D3E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FDD24890EA0D417F650FB21D5A4C37C6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"9A1562B41DFC09AF6C55ECD14D3E";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FDD24890EA0D417F650FB21D5A4C37C6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1006 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"9A1562B41DFC09AF6C55ECD14D3E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"780E97987676986969BB6996200990CA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"9A1562B41DFC09AF6C55ECD14D3E";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"780E97987676986969BB6996200990CA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1007 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"9A1562B41DFC09AF6C55ECD14D3E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C88FCCC5DD75DEEE519D28F029A2D814") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"9A1562B41DFC09AF6C55ECD14D3E";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C88FCCC5DD75DEEE519D28F029A2D814") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1008 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"9A1562B41DFC09AF6C55ECD14D3E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7689F410EEA51CEEA9E04F6210E553FE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"9A1562B41DFC09AF6C55ECD14D3E";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7689F410EEA51CEEA9E04F6210E553FE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1009 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"9A1562B41DFC09AF6C55ECD14D3E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4927007A25A542C50F47FC8B4D477D43") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"9A1562B41DFC09AF6C55ECD14D3E";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4927007A25A542C50F47FC8B4D477D43") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1010 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"9A1562B41DFC09AF6C55ECD14D3E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D150785005B519377359EA5596C90E93") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"9A1562B41DFC09AF6C55ECD14D3E";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D150785005B519377359EA5596C90E93") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1011 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"9A1562B41DFC09AF6C55ECD14D3E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AD669965E10BD2986E2BFDC288BADB24") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"9A1562B41DFC09AF6C55ECD14D3E";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AD669965E10BD2986E2BFDC288BADB24") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1012 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"9A1562B41DFC09AF6C55ECD14D3E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AD86C9BEF9AFE79C5F30BF2100C11D76") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"9A1562B41DFC09AF6C55ECD14D3E";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AD86C9BEF9AFE79C5F30BF2100C11D76") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1013 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"9A1562B41DFC09AF6C55ECD14D3E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7E7F58684DA9BCEE75720731E24DD5F9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"9A1562B41DFC09AF6C55ECD14D3E";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7E7F58684DA9BCEE75720731E24DD5F9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1014 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"9A1562B41DFC09AF6C55ECD14D3E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B86A58724DE65C8DDDEDB153E3D1E27B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"9A1562B41DFC09AF6C55ECD14D3E";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B86A58724DE65C8DDDEDB153E3D1E27B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1015 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"9A1562B41DFC09AF6C55ECD14D3E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3E73009EF0906A963E379EF7C4CADCED") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"9A1562B41DFC09AF6C55ECD14D3E";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3E73009EF0906A963E379EF7C4CADCED") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1016 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"9A1562B41DFC09AF6C55ECD14D3E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9508D499F8E92DED8B7B96F8E8C67A9D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"9A1562B41DFC09AF6C55ECD14D3E";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9508D499F8E92DED8B7B96F8E8C67A9D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1017 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"9A1562B41DFC09AF6C55ECD14D3E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8C6CCA68F99CF63D2FE1CA82962111DD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"9A1562B41DFC09AF6C55ECD14D3E";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8C6CCA68F99CF63D2FE1CA82962111DD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1018 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"9A1562B41DFC09AF6C55ECD14D3E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"39BC30A9F7488EFB1F84B3DECAA236EE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"9A1562B41DFC09AF6C55ECD14D3E";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"39BC30A9F7488EFB1F84B3DECAA236EE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1019 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"9A1562B41DFC09AF6C55ECD14D3E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F7C247132B0C1B251925DD12E98505AC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"9A1562B41DFC09AF6C55ECD14D3E";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F7C247132B0C1B251925DD12E98505AC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1020 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"9A1562B41DFC09AF6C55ECD14D3E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4D390D2661AF49837ADCE44ABC64DEA7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"9A1562B41DFC09AF6C55ECD14D3E";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4D390D2661AF49837ADCE44ABC64DEA7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1021 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"9A1562B41DFC09AF6C55ECD14D3E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EE82766D98DE8AF9AB3FC391DC50ADA2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"9A1562B41DFC09AF6C55ECD14D3E";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EE82766D98DE8AF9AB3FC391DC50ADA2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1022 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"9A1562B41DFC09AF6C55ECD14D3E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B633069E7461082CDAB5F249A89AD9C9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"9A1562B41DFC09AF6C55ECD14D3E";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B633069E7461082CDAB5F249A89AD9C9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1023 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"9A1562B41DFC09AF6C55ECD14D3E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"88FEB30DFE4BE149CA14065FF0919946") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"9A1562B41DFC09AF6C55ECD14D3E";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"88FEB30DFE4BE149CA14065FF0919946") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1024 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"9A1562B41DFC09AF6C55ECD14D3E02") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5D500028D0FB4F9CC38937707DB1F2E8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"9A1562B41DFC09AF6C55ECD14D3E02";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5D500028D0FB4F9CC38937707DB1F2E8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1025 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"9A1562B41DFC09AF6C55ECD14D3E02") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"83BE802D9D2B3CA5FEC9DA098D964871") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"9A1562B41DFC09AF6C55ECD14D3E02";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"83BE802D9D2B3CA5FEC9DA098D964871") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1026 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"9A1562B41DFC09AF6C55ECD14D3E02") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A2964603F8D97001477E035909CE29AE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"9A1562B41DFC09AF6C55ECD14D3E02";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A2964603F8D97001477E035909CE29AE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1027 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"9A1562B41DFC09AF6C55ECD14D3E02") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0601B7F940284D7D6ACC7A5AF86FF531") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"9A1562B41DFC09AF6C55ECD14D3E02";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0601B7F940284D7D6ACC7A5AF86FF531") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1028 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"9A1562B41DFC09AF6C55ECD14D3E02") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0E8746C6A53C1DEF2B4B6A4DDB2B8802") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"9A1562B41DFC09AF6C55ECD14D3E02";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0E8746C6A53C1DEF2B4B6A4DDB2B8802") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1029 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"9A1562B41DFC09AF6C55ECD14D3E02") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1A140A4AE219EFC352549125335DD2A8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"9A1562B41DFC09AF6C55ECD14D3E02";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1A140A4AE219EFC352549125335DD2A8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1030 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"9A1562B41DFC09AF6C55ECD14D3E02") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2E691BA99DC688C7E07C942060183AFA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"9A1562B41DFC09AF6C55ECD14D3E02";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2E691BA99DC688C7E07C942060183AFA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1031 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"9A1562B41DFC09AF6C55ECD14D3E02") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"13EF6A41870228A703BA46D78C90E76A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"9A1562B41DFC09AF6C55ECD14D3E02";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"13EF6A41870228A703BA46D78C90E76A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1032 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"9A1562B41DFC09AF6C55ECD14D3E02") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3E1D8BC77D601937063EA1356D6142A4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"9A1562B41DFC09AF6C55ECD14D3E02";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3E1D8BC77D601937063EA1356D6142A4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1033 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"9A1562B41DFC09AF6C55ECD14D3E02") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0F6E4E5D82FFEDAFA28A66A06BC4A1E4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"9A1562B41DFC09AF6C55ECD14D3E02";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0F6E4E5D82FFEDAFA28A66A06BC4A1E4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1034 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"9A1562B41DFC09AF6C55ECD14D3E02") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FCF22FAA907369F102CE09F048429EEB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"9A1562B41DFC09AF6C55ECD14D3E02";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FCF22FAA907369F102CE09F048429EEB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1035 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"9A1562B41DFC09AF6C55ECD14D3E02") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C7EEC463BF841EB7EE66A78E7062CC5F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"9A1562B41DFC09AF6C55ECD14D3E02";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C7EEC463BF841EB7EE66A78E7062CC5F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1036 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"9A1562B41DFC09AF6C55ECD14D3E02") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3C3F8BFBB0C903C035E2E168D54F19B3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"9A1562B41DFC09AF6C55ECD14D3E02";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3C3F8BFBB0C903C035E2E168D54F19B3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1037 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"9A1562B41DFC09AF6C55ECD14D3E02") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B65362425A3313BAF368EDF345F54C2C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"9A1562B41DFC09AF6C55ECD14D3E02";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B65362425A3313BAF368EDF345F54C2C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1038 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"9A1562B41DFC09AF6C55ECD14D3E02") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8789374A5A825C1D1BF8F22E945EE8AA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"9A1562B41DFC09AF6C55ECD14D3E02";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8789374A5A825C1D1BF8F22E945EE8AA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1039 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"9A1562B41DFC09AF6C55ECD14D3E02") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0255E842C6F9850B174C29A5EE1B4FA6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"9A1562B41DFC09AF6C55ECD14D3E02";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0255E842C6F9850B174C29A5EE1B4FA6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1040 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"9A1562B41DFC09AF6C55ECD14D3E02") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B2D4B31F6DFAC38C2F6A68C3E7B00778") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"9A1562B41DFC09AF6C55ECD14D3E02";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B2D4B31F6DFAC38C2F6A68C3E7B00778") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1041 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"9A1562B41DFC09AF6C55ECD14D3E02") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0CD28BCA5E2A018CD7170F51DEF78C92") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"9A1562B41DFC09AF6C55ECD14D3E02";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0CD28BCA5E2A018CD7170F51DEF78C92") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1042 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"9A1562B41DFC09AF6C55ECD14D3E02") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"337C7FA0952A5FA771B0BCB88355A22F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"9A1562B41DFC09AF6C55ECD14D3E02";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"337C7FA0952A5FA771B0BCB88355A22F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1043 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"9A1562B41DFC09AF6C55ECD14D3E02") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AB0B078AB53A04550DAEAA6658DBD1FF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"9A1562B41DFC09AF6C55ECD14D3E02";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AB0B078AB53A04550DAEAA6658DBD1FF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1044 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"9A1562B41DFC09AF6C55ECD14D3E02") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D73DE6BF5184CFFA10DCBDF146A80448") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"9A1562B41DFC09AF6C55ECD14D3E02";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D73DE6BF5184CFFA10DCBDF146A80448") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1045 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"9A1562B41DFC09AF6C55ECD14D3E02") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D7DDB6644920FAFE21C7FF12CED3C21A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"9A1562B41DFC09AF6C55ECD14D3E02";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D7DDB6644920FAFE21C7FF12CED3C21A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1046 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"9A1562B41DFC09AF6C55ECD14D3E02") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"042427B2FD26A18C0B8547022C5F0A95") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"9A1562B41DFC09AF6C55ECD14D3E02";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"042427B2FD26A18C0B8547022C5F0A95") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1047 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"9A1562B41DFC09AF6C55ECD14D3E02") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C23127A8FD6941EFA31AF1602DC33D17") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"9A1562B41DFC09AF6C55ECD14D3E02";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C23127A8FD6941EFA31AF1602DC33D17") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1048 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"9A1562B41DFC09AF6C55ECD14D3E02") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"44287F44401F77F440C0DEC40AD80381") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"9A1562B41DFC09AF6C55ECD14D3E02";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"44287F44401F77F440C0DEC40AD80381") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1049 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"9A1562B41DFC09AF6C55ECD14D3E02") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EF53AB434866308FF58CD6CB26D4A5F1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"9A1562B41DFC09AF6C55ECD14D3E02";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EF53AB434866308FF58CD6CB26D4A5F1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1050 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"9A1562B41DFC09AF6C55ECD14D3E02") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F637B5B24913EB5F51168AB15833CEB1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"9A1562B41DFC09AF6C55ECD14D3E02";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F637B5B24913EB5F51168AB15833CEB1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1051 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"9A1562B41DFC09AF6C55ECD14D3E02") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"43E74F7347C793996173F3ED04B0E982") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"9A1562B41DFC09AF6C55ECD14D3E02";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"43E74F7347C793996173F3ED04B0E982") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1052 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"9A1562B41DFC09AF6C55ECD14D3E02") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8D9938C99B83064767D29D212797DAC0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"9A1562B41DFC09AF6C55ECD14D3E02";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8D9938C99B83064767D29D212797DAC0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1053 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"9A1562B41DFC09AF6C55ECD14D3E02") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"376272FCD12054E1042BA479727601CB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"9A1562B41DFC09AF6C55ECD14D3E02";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"376272FCD12054E1042BA479727601CB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1054 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"9A1562B41DFC09AF6C55ECD14D3E02") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"94D909B72851979BD5C883A2124272CE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"9A1562B41DFC09AF6C55ECD14D3E02";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"94D909B72851979BD5C883A2124272CE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1055 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"9A1562B41DFC09AF6C55ECD14D3E02") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CC687944C4EE154EA442B27A668806A5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"9A1562B41DFC09AF6C55ECD14D3E02";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CC687944C4EE154EA442B27A668806A5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1056 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"9A1562B41DFC09AF6C55ECD14D3E02") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F2A5CCD74EC4FC2BB4E3466C3E83462A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"9A1562B41DFC09AF6C55ECD14D3E02";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F2A5CCD74EC4FC2BB4E3466C3E83462A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1057 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"67EF4064A3ED5F36CC0BA74D19273635") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9B074C23991F13AD9FC3B06AAC56AA8B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"67EF4064A3ED5F36CC0BA74D19273635";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9B074C23991F13AD9FC3B06AAC56AA8B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1058 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"67EF4064A3ED5F36CC0BA74D19273635") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"45E9CC26D4CF6094A2835D135C711012") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"67EF4064A3ED5F36CC0BA74D19273635";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"45E9CC26D4CF6094A2835D135C711012") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1059 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"67EF4064A3ED5F36CC0BA74D19273635") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"64C10A08B13D2C301B348443D82971CD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"67EF4064A3ED5F36CC0BA74D19273635";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"64C10A08B13D2C301B348443D82971CD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1060 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"67EF4064A3ED5F36CC0BA74D19273635") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C056FBF209CC114C3686FD402988AD52") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"67EF4064A3ED5F36CC0BA74D19273635";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C056FBF209CC114C3686FD402988AD52") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1061 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"67EF4064A3ED5F36CC0BA74D19273635") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C8D00ACDECD841DE7701ED570ACCD061") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"67EF4064A3ED5F36CC0BA74D19273635";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C8D00ACDECD841DE7701ED570ACCD061") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1062 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"67EF4064A3ED5F36CC0BA74D19273635") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DC434641ABFDB3F20E1E163FE2BA8ACB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"67EF4064A3ED5F36CC0BA74D19273635";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DC434641ABFDB3F20E1E163FE2BA8ACB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1063 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"67EF4064A3ED5F36CC0BA74D19273635") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E83E57A2D422D4F6BC36133AB1FF6299") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"67EF4064A3ED5F36CC0BA74D19273635";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E83E57A2D422D4F6BC36133AB1FF6299") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1064 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"67EF4064A3ED5F36CC0BA74D19273635") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D5B8264ACEE674965FF0C1CD5D77BF09") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"67EF4064A3ED5F36CC0BA74D19273635";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D5B8264ACEE674965FF0C1CD5D77BF09") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1065 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"67EF4064A3ED5F36CC0BA74D19273635") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F84AC7CC348445065A74262FBC861AC7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"67EF4064A3ED5F36CC0BA74D19273635";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F84AC7CC348445065A74262FBC861AC7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1066 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"67EF4064A3ED5F36CC0BA74D19273635") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C9390256CB1BB19EFEC0E1BABA23F987") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"67EF4064A3ED5F36CC0BA74D19273635";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C9390256CB1BB19EFEC0E1BABA23F987") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1067 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"67EF4064A3ED5F36CC0BA74D19273635") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3AA563A1D99735C05E848EEA99A5C688") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"67EF4064A3ED5F36CC0BA74D19273635";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3AA563A1D99735C05E848EEA99A5C688") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1068 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"67EF4064A3ED5F36CC0BA74D19273635") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"01B98868F6604286B22C2094A185943C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"67EF4064A3ED5F36CC0BA74D19273635";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"01B98868F6604286B22C2094A185943C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1069 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"67EF4064A3ED5F36CC0BA74D19273635") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FA68C7F0F92D5FF169A8667204A841D0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"67EF4064A3ED5F36CC0BA74D19273635";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FA68C7F0F92D5FF169A8667204A841D0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1070 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"67EF4064A3ED5F36CC0BA74D19273635") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"70042E4913D74F8BAF226AE99412144F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"67EF4064A3ED5F36CC0BA74D19273635";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"70042E4913D74F8BAF226AE99412144F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1071 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"67EF4064A3ED5F36CC0BA74D19273635") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"41DE7B411366002C47B2753445B9B0C9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"67EF4064A3ED5F36CC0BA74D19273635";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"41DE7B411366002C47B2753445B9B0C9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1072 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"67EF4064A3ED5F36CC0BA74D19273635") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C402A4498F1DD93A4B06AEBF3FFC17C5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"67EF4064A3ED5F36CC0BA74D19273635";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C402A4498F1DD93A4B06AEBF3FFC17C5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1073 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"67EF4064A3ED5F36CC0BA74D19273635") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7483FF14241E9FBD7320EFD936575F1B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"67EF4064A3ED5F36CC0BA74D19273635";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7483FF14241E9FBD7320EFD936575F1B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1074 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"67EF4064A3ED5F36CC0BA74D19273635") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CA85C7C117CE5DBD8B5D884B0F10D4F1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"67EF4064A3ED5F36CC0BA74D19273635";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CA85C7C117CE5DBD8B5D884B0F10D4F1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1075 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"67EF4064A3ED5F36CC0BA74D19273635") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F52B33ABDCCE03962DFA3BA252B2FA4C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"67EF4064A3ED5F36CC0BA74D19273635";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F52B33ABDCCE03962DFA3BA252B2FA4C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1076 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"67EF4064A3ED5F36CC0BA74D19273635") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6D5C4B81FCDE586451E42D7C893C899C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"67EF4064A3ED5F36CC0BA74D19273635";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6D5C4B81FCDE586451E42D7C893C899C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1077 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"67EF4064A3ED5F36CC0BA74D19273635") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"116AAAB4186093CB4C963AEB974F5C2B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"67EF4064A3ED5F36CC0BA74D19273635";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"116AAAB4186093CB4C963AEB974F5C2B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1078 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"67EF4064A3ED5F36CC0BA74D19273635") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"118AFA6F00C4A6CF7D8D78081F349A79") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"67EF4064A3ED5F36CC0BA74D19273635";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"118AFA6F00C4A6CF7D8D78081F349A79") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1079 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"67EF4064A3ED5F36CC0BA74D19273635") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C2736BB9B4C2FDBD57CFC018FDB852F6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"67EF4064A3ED5F36CC0BA74D19273635";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C2736BB9B4C2FDBD57CFC018FDB852F6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1080 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"67EF4064A3ED5F36CC0BA74D19273635") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"04666BA3B48D1DDEFF50767AFC246574") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"67EF4064A3ED5F36CC0BA74D19273635";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"04666BA3B48D1DDEFF50767AFC246574") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1081 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"67EF4064A3ED5F36CC0BA74D19273635") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"827F334F09FB2BC51C8A59DEDB3F5BE2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"67EF4064A3ED5F36CC0BA74D19273635";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"827F334F09FB2BC51C8A59DEDB3F5BE2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1082 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"67EF4064A3ED5F36CC0BA74D19273635") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2904E74801826CBEA9C651D1F733FD92") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"67EF4064A3ED5F36CC0BA74D19273635";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2904E74801826CBEA9C651D1F733FD92") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1083 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"67EF4064A3ED5F36CC0BA74D19273635") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3060F9B900F7B76E0D5C0DAB89D496D2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"67EF4064A3ED5F36CC0BA74D19273635";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3060F9B900F7B76E0D5C0DAB89D496D2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1084 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"67EF4064A3ED5F36CC0BA74D19273635") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"85B003780E23CFA83D3974F7D557B1E1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"67EF4064A3ED5F36CC0BA74D19273635";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"85B003780E23CFA83D3974F7D557B1E1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1085 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"67EF4064A3ED5F36CC0BA74D19273635") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4BCE74C2D2675A763B981A3BF67082A3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"67EF4064A3ED5F36CC0BA74D19273635";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4BCE74C2D2675A763B981A3BF67082A3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1086 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"67EF4064A3ED5F36CC0BA74D19273635") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F1353EF798C408D058612363A39159A8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"67EF4064A3ED5F36CC0BA74D19273635";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F1353EF798C408D058612363A39159A8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1087 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"67EF4064A3ED5F36CC0BA74D19273635") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"528E45BC61B5CBAA898204B8C3A52AAD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"67EF4064A3ED5F36CC0BA74D19273635";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"528E45BC61B5CBAA898204B8C3A52AAD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1088 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"67EF4064A3ED5F36CC0BA74D19273635") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0A3F354F8D0A497FF8083560B76F5EC6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"67EF4064A3ED5F36CC0BA74D19273635";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0A3F354F8D0A497FF8083560B76F5EC6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1089 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"241F0DAC2C5DDA488F0E68CADBF2CC9F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"67EF4064A3ED5F36CC0BA74D19273635") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"34F280DC0720A01AE8A9C176EF641E49") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"241F0DAC2C5DDA488F0E68CADBF2CC9F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"67EF4064A3ED5F36CC0BA74D19273635";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"34F280DC0720A01AE8A9C176EF641E49") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      wait;
   end process;

END;
