--
-- SKINNY-AEAD Reference Hardware Implementation
-- 
-- Copyright 2019:
--     Amir Moradi & Pascal Sasdrich for the SKINNY Team
--     https://sites.google.com/site/skinnycipher/
-- 
-- This program is free software; you can redistribute it and/or
-- modify it under the terms of the GNU General Public License as
-- published by the Free Software Foundation; either version 2 of the
-- License, or (at your option) any later version.
-- 
-- This program is distributed in the hope that it will be useful, but
-- WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE. See the GNU
-- General Public License for more details.
-- 

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE IEEE.std_logic_textio.all;
USE ieee.numeric_std.ALL;
USE ieee.math_real.ALL; 

ENTITY SKINNY_tk3_AEAD_encdec_M3_Test_Part1 IS
END SKINNY_tk3_AEAD_encdec_M3_Test_Part1;
 
ARCHITECTURE behavior OF SKINNY_tk3_AEAD_encdec_M3_Test_Part1 IS 
 
	constant	nl		 : integer := 0; -- 128-bit nonce
	constant	tl		 : integer := 1; --  64-bit tag     -> M3
 
 
   COMPONENT SKINNY_tk3_AEAD
	Generic (
		nl				 : integer;  -- 0: 128-bit nonce, 1: 96-bit nonce
		tl				 : integer); -- 0: 128-bit tag,   1: 64-bit tag
	Port (  
		clk          : in  STD_LOGIC;
		rst      	 : in  STD_LOGIC;
		a_data       : in  STD_LOGIC;
		enc          : in  STD_LOGIC;
		dec          : in  STD_LOGIC;
		gen_tag      : in  std_logic;
		Input1       : in  STD_LOGIC_VECTOR (127       downto 0);  -- Message or Associated Data (share 1)
		Input2       : in  STD_LOGIC_VECTOR (127       downto 0);  -- Message or Associated Data (share 2)
		N            : in  STD_LOGIC_VECTOR (127-nl*32 downto 0);
		K1           : in  STD_LOGIC_VECTOR (127       downto 0); -- Key (share 1)
		K2           : in  STD_LOGIC_VECTOR (127       downto 0); -- Key (share 2)
		Block_Size	 : in  STD_LOGIC_VECTOR (  3       downto 0); -- Size of the given block as Input (in BYTES) - 1
		Output1      : out STD_LOGIC_VECTOR (127       downto 0); -- Ciphertext (share 1)
		Output2      : out STD_LOGIC_VECTOR (127       downto 0); -- Ciphertext (share 2) 
		Tag1			 : out STD_LOGIC_VECTOR (127-tl*64 downto 0); -- Tag (share 1)
		Tag2			 : out STD_LOGIC_VECTOR (127-tl*64 downto 0); -- Tag (share 2)
		done         : out STD_LOGIC);
	END COMPONENT;
    

   --Inputs
   signal clk 			: std_logic := '0';
   signal rst 			: std_logic := '0';
   signal a_data 		: std_logic := '0';
   signal enc 			: std_logic := '0';
   signal dec 			: std_logic := '0';
   signal gen_tag 	: std_logic := '0';
   signal Input1 		: std_logic_vector(127       downto 0) := (others => '0');
   signal Input2 		: std_logic_vector(127       downto 0) := (others => '0');
   signal N 			: std_logic_vector(127-nl*32 downto 0) := (others => '0');
   signal K1 			: std_logic_vector(127       downto 0) := (others => '0');
   signal K2 			: std_logic_vector(127       downto 0) := (others => '0');
   signal Block_Size : std_logic_vector(  3       downto 0) := (others => '0');

 	--Outputs
   signal Output1		: std_logic_vector(127 downto 0);
   signal Output2		: std_logic_vector(127 downto 0);
   signal Tag1		   : std_logic_vector(127-tl*64 downto 0);
   signal Tag2		   : std_logic_vector(127-tl*64 downto 0);
   signal done 		: std_logic;

   signal Input 		: std_logic_vector(127 downto 0) := (others => '0');
   signal K 			: std_logic_vector(127 downto 0) := (others => '0');
   signal Output		: std_logic_vector(127 downto 0);
   signal Tag		   : std_logic_vector(127-tl*64 downto 0);

	signal Mask1		: std_logic_vector(127 downto 0);
	signal Mask2		: std_logic_vector(127 downto 0);
	

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
 	type INT_ARRAY  is array (integer range <>) of integer range 0 to 255;
	type REAL_ARRAY is array (integer range <>) of real;
	type BYTE_ARRAY is array (integer range <>) of std_logic_vector(7 downto 0);

	signal r: INT_ARRAY (31 downto 0);
	signal m: BYTE_ARRAY(31 downto 0);

BEGIN
 
  	maskgen: process
		 variable seed1, seed2: positive;        -- seed values for random generator
		 variable rand: REAL_ARRAY(31 downto 0); -- random real-number value in range 0 to 1.0  
		 variable range_of_rand : real := 256.0; -- the range of random values created will be 0 to +255.
	begin
		 
		FOR i in 0 to 31 loop
			uniform(seed1, seed2, rand(i));   -- generate random number
			r(i) <= integer(TRUNC(rand(i)*range_of_rand));  -- rescale to 0...255, convert integer part 
			m(i) <= std_logic_vector(to_unsigned(r(i), m(i)'length));
		end loop;
		
		wait for clk_period;
	end process;  

	---------
	
	maskassign: FOR i in 0 to 15 GENERATE
		Mask1(i*8+7 downto i*8)	<= m(i);
		Mask2(i*8+7 downto i*8)	<= m(16+i);
	END GENERATE;

	---------
 
   uut: SKINNY_tk3_AEAD 
	GENERIC MAP (
		nl		=> nl,
		tl		=> tl)
	PORT MAP (
		clk 			=> clk,
		rst 			=> rst,
		a_data 		=> a_data,
		enc 			=> enc,
		dec			=> dec,
		gen_tag 		=> gen_tag,
		Input1 		=> Input1,
		Input2 		=> Input2,
		N 				=> N,
		K1				=> K1,
		K2				=> K2,
		Block_Size 	=> Block_Size,
		Output1 		=> Output1,
		Output2 		=> Output2,
		Tag1			=> Tag1,
		Tag2			=> Tag2,
		done 			=> done);

	Input1	<= Input XOR Mask1;
	Input2	<= Mask1;

	K1			<= K XOR Mask2;
	K2			<= Mask2;

	Output	<= Output1 XOR Output2;
	Tag		<= Tag1 XOR Tag2;

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      --------- test no. 1 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"62B08C0557EDCC94") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 2 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"ECCD324D36BFF667") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 3 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BF80E07AF4D1916F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 4 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"165482D6E01D234E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 5 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A8741920DA4B04ED") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 6 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0752C75717EB3A96") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 7 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B530CAA5A9C69486") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 8 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DEA9A081C5DBF74B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 9 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"044F82139B4FB39D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 10 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AB47BB9205EEA704") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 11 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0DBEEA9A2FD2252E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 12 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B4B4DA869FA9C73A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 13 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D4FAA611D313E648") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 14 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FC5540B1CFD8E4E0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 15 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"872D62831CF0C36B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 16 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0AAB4B55C8A1B1BF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 17 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E414ED04167F946B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 18 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C384F572382054C3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 19 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EFEA7517D1CE3292") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 20 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"50239F30A567BCD0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 21 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BDF27F4D7D2F9581") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 22 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"99217CEC6E294D18") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 23 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EC03FD0F5ECA21EC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 24 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"90DFCCC23FB814B8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 25 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2EFDCC8CBA4A15BD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 26 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BCEA51A38385C4EB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 27 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"716D84F17AA2BBA2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 28 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D6F14EC029B71B8C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 29 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3CD780C215026F8D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 30 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6405E297CAC12A56") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 31 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7EC61B0F6A28B310") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 32 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"69217A69416D623E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 33 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6BFA0110F0335845") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 34 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"80") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D922B9DBC87717CF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"80";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D922B9DBC87717CF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 35 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"80") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"575F0793A9252D3C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"80";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"575F0793A9252D3C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 36 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"80") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0412D5A46B4B4A34") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"80";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0412D5A46B4B4A34") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 37 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"80") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"ADC6B7087F87F815") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"80";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"ADC6B7087F87F815") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 38 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"80") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"13E62CFE45D1DFB6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"80";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"13E62CFE45D1DFB6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 39 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"80") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BCC0F2898871E1CD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"80";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BCC0F2898871E1CD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 40 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"80") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0EA2FF7B365C4FDD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"80";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0EA2FF7B365C4FDD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 41 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"80") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"653B955F5A412C10") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"80";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"653B955F5A412C10") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 42 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"80") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BFDDB7CD04D568C6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"80";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BFDDB7CD04D568C6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 43 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"80") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"10D58E4C9A747C5F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"80";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"10D58E4C9A747C5F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 44 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"80") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B62CDF44B048FE75") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"80";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B62CDF44B048FE75") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 45 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"80") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0F26EF5800331C61") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"80";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0F26EF5800331C61") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 46 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"80") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6F6893CF4C893D13") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"80";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6F6893CF4C893D13") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 47 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"80") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"47C7756F50423FBB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"80";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"47C7756F50423FBB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 48 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"80") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3CBF575D836A1830") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"80";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3CBF575D836A1830") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 49 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"80") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B1397E8B573B6AE4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"80";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B1397E8B573B6AE4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 50 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"80") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5F86D8DA89E54F30") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"80";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5F86D8DA89E54F30") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 51 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"80") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7816C0ACA7BA8F98") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"80";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7816C0ACA7BA8F98") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 52 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"80") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"547840C94E54E9C9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"80";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"547840C94E54E9C9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 53 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"80") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EBB1AAEE3AFD678B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"80";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EBB1AAEE3AFD678B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 54 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"80") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"06604A93E2B54EDA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"80";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"06604A93E2B54EDA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 55 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"80") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"22B34932F1B39643") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"80";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"22B34932F1B39643") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 56 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"80") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5791C8D1C150FAB7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"80";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5791C8D1C150FAB7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 57 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"80") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2B4DF91CA022CFE3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"80";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2B4DF91CA022CFE3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 58 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"80") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"956FF95225D0CEE6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"80";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"956FF95225D0CEE6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 59 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"80") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0778647D1C1F1FB0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"80";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0778647D1C1F1FB0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 60 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"80") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CAFFB12FE53860F9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"80";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CAFFB12FE53860F9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 61 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"80") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6D637B1EB62DC0D7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"80";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6D637B1EB62DC0D7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 62 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"80") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8745B51C8A98B4D6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"80";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8745B51C8A98B4D6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 63 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"80") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DF97D749555BF10D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"80";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DF97D749555BF10D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 64 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"80") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C5542ED1F5B2684B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"80";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C5542ED1F5B2684B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 65 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"80") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D2B34FB7DEF7B965") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"80";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D2B34FB7DEF7B965") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 66 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"80") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D06834CE6FA9831E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"80";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"00") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D06834CE6FA9831E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 67 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"80E4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B10164FB19931A67") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"80E4";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B10164FB19931A67") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 68 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"80E4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3F7CDAB378C12094") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"80E4";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3F7CDAB378C12094") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 69 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"80E4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6C310884BAAF479C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"80E4";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6C310884BAAF479C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 70 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"80E4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C5E56A28AE63F5BD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"80E4";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C5E56A28AE63F5BD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 71 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"80E4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7BC5F1DE9435D21E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"80E4";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7BC5F1DE9435D21E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 72 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"80E4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D4E32FA95995EC65") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"80E4";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D4E32FA95995EC65") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 73 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"80E4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6681225BE7B84275") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"80E4";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6681225BE7B84275") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 74 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"80E4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0D18487F8BA521B8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"80E4";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0D18487F8BA521B8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 75 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"80E4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D7FE6AEDD531656E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"80E4";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D7FE6AEDD531656E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 76 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"80E4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"78F6536C4B9071F7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"80E4";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"78F6536C4B9071F7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 77 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"80E4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DE0F026461ACF3DD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"80E4";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DE0F026461ACF3DD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 78 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"80E4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"67053278D1D711C9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"80E4";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"67053278D1D711C9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 79 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"80E4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"074B4EEF9D6D30BB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"80E4";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"074B4EEF9D6D30BB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 80 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"80E4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2FE4A84F81A63213") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"80E4";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2FE4A84F81A63213") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 81 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"80E4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"549C8A7D528E1598") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"80E4";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"549C8A7D528E1598") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 82 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"80E4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D91AA3AB86DF674C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"80E4";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D91AA3AB86DF674C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 83 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"80E4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"37A505FA58014298") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"80E4";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"37A505FA58014298") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 84 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"80E4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"10351D8C765E8230") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"80E4";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"10351D8C765E8230") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 85 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"80E4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3C5B9DE99FB0E461") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"80E4";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3C5B9DE99FB0E461") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 86 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"80E4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"839277CEEB196A23") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"80E4";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"839277CEEB196A23") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 87 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"80E4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6E4397B333514372") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"80E4";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6E4397B333514372") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 88 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"80E4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4A90941220579BEB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"80E4";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4A90941220579BEB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 89 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"80E4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3FB215F110B4F71F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"80E4";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3FB215F110B4F71F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 90 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"80E4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"436E243C71C6C24B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"80E4";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"436E243C71C6C24B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 91 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"80E4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FD4C2472F434C34E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"80E4";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FD4C2472F434C34E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 92 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"80E4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6F5BB95DCDFB1218") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"80E4";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6F5BB95DCDFB1218") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 93 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"80E4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A2DC6C0F34DC6D51") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"80E4";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A2DC6C0F34DC6D51") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 94 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"80E4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0540A63E67C9CD7F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"80E4";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0540A63E67C9CD7F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 95 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"80E4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EF66683C5B7CB97E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"80E4";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EF66683C5B7CB97E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 96 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"80E4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B7B40A6984BFFCA5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"80E4";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B7B40A6984BFFCA5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 97 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"80E4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AD77F3F1245665E3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"80E4";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AD77F3F1245665E3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 98 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"80E4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BA9092970F13B4CD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"80E4";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BA9092970F13B4CD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 99 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"80E4") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B84BE9EEBE4D8EB6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"80E4";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"0001") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B84BE9EEBE4D8EB6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 100 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"80E435") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A8357BAACAEA1CCB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"80E435";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A8357BAACAEA1CCB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 101 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"80E435") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2648C5E2ABB82638") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"80E435";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2648C5E2ABB82638") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 102 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"80E435") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"750517D569D64130") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"80E435";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"750517D569D64130") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 103 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"80E435") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DCD175797D1AF311") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"80E435";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DCD175797D1AF311") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 104 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"80E435") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"62F1EE8F474CD4B2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"80E435";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"62F1EE8F474CD4B2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 105 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"80E435") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CDD730F88AECEAC9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"80E435";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CDD730F88AECEAC9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 106 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"80E435") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7FB53D0A34C144D9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"80E435";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7FB53D0A34C144D9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 107 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"80E435") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"142C572E58DC2714") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"80E435";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"142C572E58DC2714") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 108 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"80E435") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CECA75BC064863C2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"80E435";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CECA75BC064863C2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 109 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"80E435") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"61C24C3D98E9775B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"80E435";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"61C24C3D98E9775B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 110 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"80E435") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C73B1D35B2D5F571") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"80E435";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C73B1D35B2D5F571") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 111 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"80E435") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7E312D2902AE1765") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"80E435";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7E312D2902AE1765") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 112 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"80E435") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1E7F51BE4E143617") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"80E435";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1E7F51BE4E143617") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 113 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"80E435") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"36D0B71E52DF34BF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"80E435";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"36D0B71E52DF34BF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 114 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"80E435") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4DA8952C81F71334") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"80E435";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4DA8952C81F71334") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 115 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"80E435") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C02EBCFA55A661E0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"80E435";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C02EBCFA55A661E0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 116 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"80E435") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2E911AAB8B784434") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"80E435";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2E911AAB8B784434") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 117 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"80E435") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"090102DDA527849C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"80E435";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"090102DDA527849C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 118 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"80E435") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"256F82B84CC9E2CD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"80E435";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"256F82B84CC9E2CD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 119 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"80E435") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9AA6689F38606C8F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"80E435";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9AA6689F38606C8F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 120 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"80E435") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"777788E2E02845DE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"80E435";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"777788E2E02845DE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 121 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"80E435") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"53A48B43F32E9D47") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"80E435";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"53A48B43F32E9D47") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 122 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"80E435") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"26860AA0C3CDF1B3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"80E435";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"26860AA0C3CDF1B3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 123 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"80E435") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5A5A3B6DA2BFC4E7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"80E435";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5A5A3B6DA2BFC4E7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 124 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"80E435") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E4783B23274DC5E2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"80E435";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E4783B23274DC5E2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 125 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"80E435") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"766FA60C1E8214B4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"80E435";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"766FA60C1E8214B4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 126 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"80E435") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BBE8735EE7A56BFD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"80E435";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BBE8735EE7A56BFD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 127 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"80E435") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1C74B96FB4B0CBD3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"80E435";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1C74B96FB4B0CBD3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 128 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"80E435") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F652776D8805BFD2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"80E435";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F652776D8805BFD2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 129 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"80E435") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AE80153857C6FA09") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"80E435";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AE80153857C6FA09") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 130 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"80E435") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B443ECA0F72F634F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"80E435";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B443ECA0F72F634F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 131 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"80E435") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A3A48DC6DC6AB261") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"80E435";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A3A48DC6DC6AB261") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 132 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"80E435") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A17FF6BF6D34881A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"80E435";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"000102") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A17FF6BF6D34881A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 133 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"80E4351A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E3C0D6F40A3D756E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"80E4351A";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E3C0D6F40A3D756E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 134 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"80E4351A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6DBD68BC6B6F4F9D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"80E4351A";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6DBD68BC6B6F4F9D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 135 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"80E4351A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3EF0BA8BA9012895") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"80E4351A";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3EF0BA8BA9012895") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 136 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"80E4351A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9724D827BDCD9AB4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"80E4351A";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9724D827BDCD9AB4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 137 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"80E4351A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"290443D1879BBD17") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"80E4351A";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"290443D1879BBD17") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 138 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"80E4351A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"86229DA64A3B836C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"80E4351A";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"86229DA64A3B836C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 139 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"80E4351A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"34409054F4162D7C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"80E4351A";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"34409054F4162D7C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 140 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"80E4351A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5FD9FA70980B4EB1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"80E4351A";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5FD9FA70980B4EB1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 141 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"80E4351A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"853FD8E2C69F0A67") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"80E4351A";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"853FD8E2C69F0A67") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 142 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"80E4351A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2A37E163583E1EFE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"80E4351A";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2A37E163583E1EFE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 143 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"80E4351A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8CCEB06B72029CD4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"80E4351A";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8CCEB06B72029CD4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 144 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"80E4351A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"35C48077C2797EC0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"80E4351A";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"35C48077C2797EC0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 145 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"80E4351A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"558AFCE08EC35FB2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"80E4351A";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"558AFCE08EC35FB2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 146 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"80E4351A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7D251A4092085D1A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"80E4351A";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7D251A4092085D1A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 147 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"80E4351A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"065D387241207A91") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"80E4351A";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"065D387241207A91") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 148 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"80E4351A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8BDB11A495710845") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"80E4351A";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8BDB11A495710845") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 149 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"80E4351A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6564B7F54BAF2D91") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"80E4351A";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6564B7F54BAF2D91") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 150 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"80E4351A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"42F4AF8365F0ED39") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"80E4351A";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"42F4AF8365F0ED39") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 151 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"80E4351A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6E9A2FE68C1E8B68") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"80E4351A";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6E9A2FE68C1E8B68") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 152 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"80E4351A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D153C5C1F8B7052A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"80E4351A";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D153C5C1F8B7052A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 153 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"80E4351A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3C8225BC20FF2C7B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"80E4351A";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3C8225BC20FF2C7B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 154 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"80E4351A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1851261D33F9F4E2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"80E4351A";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1851261D33F9F4E2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 155 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"80E4351A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6D73A7FE031A9816") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"80E4351A";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6D73A7FE031A9816") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 156 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"80E4351A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"11AF96336268AD42") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"80E4351A";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"11AF96336268AD42") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 157 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"80E4351A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AF8D967DE79AAC47") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"80E4351A";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AF8D967DE79AAC47") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 158 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"80E4351A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3D9A0B52DE557D11") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"80E4351A";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3D9A0B52DE557D11") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 159 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"80E4351A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F01DDE0027720258") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"80E4351A";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F01DDE0027720258") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 160 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"80E4351A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"578114317467A276") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"80E4351A";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"578114317467A276") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 161 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"80E4351A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BDA7DA3348D2D677") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"80E4351A";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BDA7DA3348D2D677") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 162 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"80E4351A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E575B866971193AC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"80E4351A";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E575B866971193AC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 163 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"80E4351A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FFB641FE37F80AEA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"80E4351A";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FFB641FE37F80AEA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 164 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"80E4351A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E85120981CBDDBC4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"80E4351A";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E85120981CBDDBC4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 165 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"80E4351A") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EA8A5BE1ADE3E1BF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"80E4351A";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"00010203") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EA8A5BE1ADE3E1BF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 166 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"80E4351A76") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1E5D9F7B94431FCC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"80E4351A76";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1E5D9F7B94431FCC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 167 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"80E4351A76") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"90202133F511253F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"80E4351A76";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"90202133F511253F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 168 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"80E4351A76") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C36DF304377F4237") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"80E4351A76";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C36DF304377F4237") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 169 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"80E4351A76") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6AB991A823B3F016") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"80E4351A76";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6AB991A823B3F016") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 170 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"80E4351A76") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D4990A5E19E5D7B5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"80E4351A76";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D4990A5E19E5D7B5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 171 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"80E4351A76") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7BBFD429D445E9CE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"80E4351A76";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7BBFD429D445E9CE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 172 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"80E4351A76") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C9DDD9DB6A6847DE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"80E4351A76";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C9DDD9DB6A6847DE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 173 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"80E4351A76") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A244B3FF06752413") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"80E4351A76";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A244B3FF06752413") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 174 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"80E4351A76") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"78A2916D58E160C5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"80E4351A76";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"78A2916D58E160C5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 175 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"80E4351A76") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D7AAA8ECC640745C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"80E4351A76";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D7AAA8ECC640745C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 176 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"80E4351A76") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7153F9E4EC7CF676") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"80E4351A76";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7153F9E4EC7CF676") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 177 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"80E4351A76") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C859C9F85C071462") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"80E4351A76";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C859C9F85C071462") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 178 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"80E4351A76") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A817B56F10BD3510") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"80E4351A76";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A817B56F10BD3510") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 179 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"80E4351A76") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"80B853CF0C7637B8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"80E4351A76";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"80B853CF0C7637B8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 180 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"80E4351A76") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FBC071FDDF5E1033") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"80E4351A76";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FBC071FDDF5E1033") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 181 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"80E4351A76") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7646582B0B0F62E7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"80E4351A76";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7646582B0B0F62E7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 182 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"80E4351A76") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"98F9FE7AD5D14733") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"80E4351A76";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"98F9FE7AD5D14733") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 183 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"80E4351A76") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BF69E60CFB8E879B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"80E4351A76";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BF69E60CFB8E879B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 184 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"80E4351A76") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"930766691260E1CA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"80E4351A76";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"930766691260E1CA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 185 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"80E4351A76") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2CCE8C4E66C96F88") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"80E4351A76";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2CCE8C4E66C96F88") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 186 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"80E4351A76") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C11F6C33BE8146D9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"80E4351A76";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C11F6C33BE8146D9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 187 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"80E4351A76") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E5CC6F92AD879E40") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"80E4351A76";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E5CC6F92AD879E40") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 188 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"80E4351A76") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"90EEEE719D64F2B4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"80E4351A76";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"90EEEE719D64F2B4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 189 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"80E4351A76") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EC32DFBCFC16C7E0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"80E4351A76";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EC32DFBCFC16C7E0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 190 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"80E4351A76") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5210DFF279E4C6E5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"80E4351A76";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5210DFF279E4C6E5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 191 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"80E4351A76") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C00742DD402B17B3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"80E4351A76";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C00742DD402B17B3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 192 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"80E4351A76") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0D80978FB90C68FA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"80E4351A76";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0D80978FB90C68FA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 193 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"80E4351A76") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AA1C5DBEEA19C8D4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"80E4351A76";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AA1C5DBEEA19C8D4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 194 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"80E4351A76") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"403A93BCD6ACBCD5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"80E4351A76";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"403A93BCD6ACBCD5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 195 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"80E4351A76") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"18E8F1E9096FF90E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"80E4351A76";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"18E8F1E9096FF90E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 196 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"80E4351A76") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"022B0871A9866048") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"80E4351A76";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"022B0871A9866048") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 197 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"80E4351A76") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"15CC691782C3B166") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"80E4351A76";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"15CC691782C3B166") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 198 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"80E4351A76") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1717126E339D8B1D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"80E4351A76";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"0001020304") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1717126E339D8B1D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 199 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"80E4351A76EF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0E401FAD7CA70EE9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"80E4351A76EF";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0E401FAD7CA70EE9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 200 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"80E4351A76EF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"803DA1E51DF5341A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"80E4351A76EF";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"803DA1E51DF5341A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 201 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"80E4351A76EF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D37073D2DF9B5312") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"80E4351A76EF";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D37073D2DF9B5312") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 202 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"80E4351A76EF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7AA4117ECB57E133") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"80E4351A76EF";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7AA4117ECB57E133") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 203 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"80E4351A76EF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C4848A88F101C690") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"80E4351A76EF";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C4848A88F101C690") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 204 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"80E4351A76EF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6BA254FF3CA1F8EB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"80E4351A76EF";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6BA254FF3CA1F8EB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 205 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"80E4351A76EF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D9C0590D828C56FB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"80E4351A76EF";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D9C0590D828C56FB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 206 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"80E4351A76EF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B2593329EE913536") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"80E4351A76EF";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B2593329EE913536") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 207 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"80E4351A76EF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"68BF11BBB00571E0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"80E4351A76EF";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"68BF11BBB00571E0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 208 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"80E4351A76EF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C7B7283A2EA46579") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"80E4351A76EF";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C7B7283A2EA46579") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 209 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"80E4351A76EF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"614E79320498E753") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"80E4351A76EF";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"614E79320498E753") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 210 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"80E4351A76EF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D844492EB4E30547") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"80E4351A76EF";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D844492EB4E30547") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 211 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"80E4351A76EF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B80A35B9F8592435") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"80E4351A76EF";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B80A35B9F8592435") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 212 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"80E4351A76EF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"90A5D319E492269D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"80E4351A76EF";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"90A5D319E492269D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 213 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"80E4351A76EF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EBDDF12B37BA0116") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"80E4351A76EF";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EBDDF12B37BA0116") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 214 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"80E4351A76EF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"665BD8FDE3EB73C2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"80E4351A76EF";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"665BD8FDE3EB73C2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 215 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"80E4351A76EF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"88E47EAC3D355616") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"80E4351A76EF";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"88E47EAC3D355616") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 216 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"80E4351A76EF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AF7466DA136A96BE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"80E4351A76EF";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AF7466DA136A96BE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 217 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"80E4351A76EF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"831AE6BFFA84F0EF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"80E4351A76EF";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"831AE6BFFA84F0EF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 218 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"80E4351A76EF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3CD30C988E2D7EAD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"80E4351A76EF";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3CD30C988E2D7EAD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 219 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"80E4351A76EF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D102ECE5566557FC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"80E4351A76EF";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D102ECE5566557FC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 220 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"80E4351A76EF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F5D1EF4445638F65") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"80E4351A76EF";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F5D1EF4445638F65") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 221 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"80E4351A76EF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"80F36EA77580E391") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"80E4351A76EF";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"80F36EA77580E391") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 222 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"80E4351A76EF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FC2F5F6A14F2D6C5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"80E4351A76EF";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FC2F5F6A14F2D6C5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 223 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"80E4351A76EF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"420D5F249100D7C0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"80E4351A76EF";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"420D5F249100D7C0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 224 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"80E4351A76EF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D01AC20BA8CF0696") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"80E4351A76EF";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D01AC20BA8CF0696") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 225 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"80E4351A76EF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1D9D175951E879DF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"80E4351A76EF";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1D9D175951E879DF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 226 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"80E4351A76EF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BA01DD6802FDD9F1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"80E4351A76EF";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BA01DD6802FDD9F1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 227 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"80E4351A76EF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5027136A3E48ADF0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"80E4351A76EF";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5027136A3E48ADF0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 228 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"80E4351A76EF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"08F5713FE18BE82B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"80E4351A76EF";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"08F5713FE18BE82B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 229 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"80E4351A76EF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"123688A74162716D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"80E4351A76EF";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"123688A74162716D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 230 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"80E4351A76EF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"05D1E9C16A27A043") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"80E4351A76EF";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"05D1E9C16A27A043") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 231 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"80E4351A76EF") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"070A92B8DB799A38") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"80E4351A76EF";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"000102030405") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"070A92B8DB799A38") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 232 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"80E4351A76EF78") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E1F43793EBDD39AA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"80E4351A76EF78";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E1F43793EBDD39AA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 233 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"80E4351A76EF78") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6F8989DB8A8F0359") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"80E4351A76EF78";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6F8989DB8A8F0359") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 234 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"80E4351A76EF78") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3CC45BEC48E16451") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"80E4351A76EF78";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3CC45BEC48E16451") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 235 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"80E4351A76EF78") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"951039405C2DD670") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"80E4351A76EF78";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"951039405C2DD670") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 236 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"80E4351A76EF78") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2B30A2B6667BF1D3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"80E4351A76EF78";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2B30A2B6667BF1D3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 237 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"80E4351A76EF78") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"84167CC1ABDBCFA8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"80E4351A76EF78";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"84167CC1ABDBCFA8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 238 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"80E4351A76EF78") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3674713315F661B8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"80E4351A76EF78";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3674713315F661B8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 239 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"80E4351A76EF78") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5DED1B1779EB0275") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"80E4351A76EF78";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5DED1B1779EB0275") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 240 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"80E4351A76EF78") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"870B3985277F46A3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"80E4351A76EF78";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"870B3985277F46A3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 241 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"80E4351A76EF78") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"28030004B9DE523A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"80E4351A76EF78";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"28030004B9DE523A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 242 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"80E4351A76EF78") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8EFA510C93E2D010") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"80E4351A76EF78";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8EFA510C93E2D010") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 243 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"80E4351A76EF78") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"37F0611023993204") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"80E4351A76EF78";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"37F0611023993204") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 244 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"80E4351A76EF78") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"57BE1D876F231376") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"80E4351A76EF78";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"57BE1D876F231376") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 245 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"80E4351A76EF78") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7F11FB2773E811DE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"80E4351A76EF78";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7F11FB2773E811DE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 246 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"80E4351A76EF78") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0469D915A0C03655") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"80E4351A76EF78";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0469D915A0C03655") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 247 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"80E4351A76EF78") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"89EFF0C374914481") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"80E4351A76EF78";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"89EFF0C374914481") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 248 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"80E4351A76EF78") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"67505692AA4F6155") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"80E4351A76EF78";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"67505692AA4F6155") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 249 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"80E4351A76EF78") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"40C04EE48410A1FD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"80E4351A76EF78";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"40C04EE48410A1FD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 250 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"80E4351A76EF78") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6CAECE816DFEC7AC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"80E4351A76EF78";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6CAECE816DFEC7AC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 251 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"80E4351A76EF78") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D36724A6195749EE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"80E4351A76EF78";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D36724A6195749EE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 252 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"80E4351A76EF78") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3EB6C4DBC11F60BF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"80E4351A76EF78";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3EB6C4DBC11F60BF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 253 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"80E4351A76EF78") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1A65C77AD219B826") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"80E4351A76EF78";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1A65C77AD219B826") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 254 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"80E4351A76EF78") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6F474699E2FAD4D2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"80E4351A76EF78";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6F474699E2FAD4D2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 255 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"80E4351A76EF78") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"139B77548388E186") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"80E4351A76EF78";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"139B77548388E186") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 256 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"80E4351A76EF78") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"ADB9771A067AE083") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"80E4351A76EF78";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"ADB9771A067AE083") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 257 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"80E4351A76EF78") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3FAEEA353FB531D5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"80E4351A76EF78";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3FAEEA353FB531D5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 258 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"80E4351A76EF78") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F2293F67C6924E9C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"80E4351A76EF78";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F2293F67C6924E9C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 259 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"80E4351A76EF78") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"55B5F5569587EEB2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"80E4351A76EF78";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"55B5F5569587EEB2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 260 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"80E4351A76EF78") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BF933B54A9329AB3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"80E4351A76EF78";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BF933B54A9329AB3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 261 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"80E4351A76EF78") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E741590176F1DF68") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"80E4351A76EF78";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E741590176F1DF68") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 262 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"80E4351A76EF78") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FD82A099D618462E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"80E4351A76EF78";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FD82A099D618462E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 263 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"80E4351A76EF78") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EA65C1FFFD5D9700") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"80E4351A76EF78";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EA65C1FFFD5D9700") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 264 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"80E4351A76EF78") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E8BEBA864C03AD7B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"80E4351A76EF78";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"00010203040506") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E8BEBA864C03AD7B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 265 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"80E4351A76EF7818") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FD221747EEDDD4F6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"80E4351A76EF7818";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FD221747EEDDD4F6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 266 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"80E4351A76EF7818") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"735FA90F8F8FEE05") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"80E4351A76EF7818";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"735FA90F8F8FEE05") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 267 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"80E4351A76EF7818") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"20127B384DE1890D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"80E4351A76EF7818";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"20127B384DE1890D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 268 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"80E4351A76EF7818") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"89C61994592D3B2C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"80E4351A76EF7818";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"89C61994592D3B2C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 269 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"80E4351A76EF7818") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"37E68262637B1C8F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"80E4351A76EF7818";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"37E68262637B1C8F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 270 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"80E4351A76EF7818") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"98C05C15AEDB22F4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"80E4351A76EF7818";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"98C05C15AEDB22F4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 271 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"80E4351A76EF7818") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2AA251E710F68CE4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"80E4351A76EF7818";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2AA251E710F68CE4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 272 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"80E4351A76EF7818") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"413B3BC37CEBEF29") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"80E4351A76EF7818";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"413B3BC37CEBEF29") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 273 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"80E4351A76EF7818") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9BDD1951227FABFF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"80E4351A76EF7818";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9BDD1951227FABFF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 274 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"80E4351A76EF7818") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"34D520D0BCDEBF66") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"80E4351A76EF7818";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"34D520D0BCDEBF66") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 275 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"80E4351A76EF7818") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"922C71D896E23D4C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"80E4351A76EF7818";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"922C71D896E23D4C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 276 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"80E4351A76EF7818") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2B2641C42699DF58") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"80E4351A76EF7818";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2B2641C42699DF58") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 277 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"80E4351A76EF7818") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4B683D536A23FE2A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"80E4351A76EF7818";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4B683D536A23FE2A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 278 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"80E4351A76EF7818") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"63C7DBF376E8FC82") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"80E4351A76EF7818";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"63C7DBF376E8FC82") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 279 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"80E4351A76EF7818") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"18BFF9C1A5C0DB09") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"80E4351A76EF7818";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"18BFF9C1A5C0DB09") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 280 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"80E4351A76EF7818") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9539D0177191A9DD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"80E4351A76EF7818";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9539D0177191A9DD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 281 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"80E4351A76EF7818") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7B867646AF4F8C09") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"80E4351A76EF7818";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7B867646AF4F8C09") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 282 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"80E4351A76EF7818") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5C166E3081104CA1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"80E4351A76EF7818";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5C166E3081104CA1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 283 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"80E4351A76EF7818") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7078EE5568FE2AF0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"80E4351A76EF7818";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7078EE5568FE2AF0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 284 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"80E4351A76EF7818") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CFB104721C57A4B2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"80E4351A76EF7818";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CFB104721C57A4B2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 285 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"80E4351A76EF7818") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2260E40FC41F8DE3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"80E4351A76EF7818";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2260E40FC41F8DE3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 286 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"80E4351A76EF7818") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"06B3E7AED719557A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"80E4351A76EF7818";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"06B3E7AED719557A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 287 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"80E4351A76EF7818") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7391664DE7FA398E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"80E4351A76EF7818";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7391664DE7FA398E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 288 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"80E4351A76EF7818") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0F4D578086880CDA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"80E4351A76EF7818";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0F4D578086880CDA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 289 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"80E4351A76EF7818") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B16F57CE037A0DDF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"80E4351A76EF7818";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B16F57CE037A0DDF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 290 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"80E4351A76EF7818") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2378CAE13AB5DC89") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"80E4351A76EF7818";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2378CAE13AB5DC89") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 291 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"80E4351A76EF7818") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EEFF1FB3C392A3C0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"80E4351A76EF7818";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EEFF1FB3C392A3C0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 292 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"80E4351A76EF7818") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4963D582908703EE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"80E4351A76EF7818";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4963D582908703EE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 293 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"80E4351A76EF7818") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A3451B80AC3277EF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"80E4351A76EF7818";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A3451B80AC3277EF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 294 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"80E4351A76EF7818") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FB9779D573F13234") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"80E4351A76EF7818";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FB9779D573F13234") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 295 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"80E4351A76EF7818") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E154804DD318AB72") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"80E4351A76EF7818";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E154804DD318AB72") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 296 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"80E4351A76EF7818") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F6B3E12BF85D7A5C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"80E4351A76EF7818";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F6B3E12BF85D7A5C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 297 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"80E4351A76EF7818") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F4689A5249034027") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"80E4351A76EF7818";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"0001020304050607") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F4689A5249034027") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 298 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"80E4351A76EF78185D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1BE92B224F336584") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"80E4351A76EF78185D";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1BE92B224F336584") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 299 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"80E4351A76EF78185D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9594956A2E615F77") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"80E4351A76EF78185D";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9594956A2E615F77") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 300 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"80E4351A76EF78185D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C6D9475DEC0F387F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"80E4351A76EF78185D";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C6D9475DEC0F387F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 301 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"80E4351A76EF78185D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6F0D25F1F8C38A5E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"80E4351A76EF78185D";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6F0D25F1F8C38A5E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 302 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"80E4351A76EF78185D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D12DBE07C295ADFD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"80E4351A76EF78185D";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D12DBE07C295ADFD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 303 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"80E4351A76EF78185D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7E0B60700F359386") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"80E4351A76EF78185D";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7E0B60700F359386") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 304 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"80E4351A76EF78185D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CC696D82B1183D96") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"80E4351A76EF78185D";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CC696D82B1183D96") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 305 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"80E4351A76EF78185D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A7F007A6DD055E5B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"80E4351A76EF78185D";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A7F007A6DD055E5B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 306 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"80E4351A76EF78185D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7D16253483911A8D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"80E4351A76EF78185D";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7D16253483911A8D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 307 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"80E4351A76EF78185D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D21E1CB51D300E14") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"80E4351A76EF78185D";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D21E1CB51D300E14") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 308 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"80E4351A76EF78185D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"74E74DBD370C8C3E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"80E4351A76EF78185D";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"74E74DBD370C8C3E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 309 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"80E4351A76EF78185D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CDED7DA187776E2A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"80E4351A76EF78185D";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CDED7DA187776E2A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 310 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"80E4351A76EF78185D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"ADA30136CBCD4F58") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"80E4351A76EF78185D";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"ADA30136CBCD4F58") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 311 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"80E4351A76EF78185D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"850CE796D7064DF0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"80E4351A76EF78185D";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"850CE796D7064DF0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 312 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"80E4351A76EF78185D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FE74C5A4042E6A7B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"80E4351A76EF78185D";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FE74C5A4042E6A7B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 313 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"80E4351A76EF78185D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"73F2EC72D07F18AF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"80E4351A76EF78185D";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"73F2EC72D07F18AF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 314 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"80E4351A76EF78185D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9D4D4A230EA13D7B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"80E4351A76EF78185D";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9D4D4A230EA13D7B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 315 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"80E4351A76EF78185D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BADD525520FEFDD3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"80E4351A76EF78185D";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BADD525520FEFDD3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 316 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"80E4351A76EF78185D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"96B3D230C9109B82") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"80E4351A76EF78185D";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"96B3D230C9109B82") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 317 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"80E4351A76EF78185D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"297A3817BDB915C0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"80E4351A76EF78185D";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"297A3817BDB915C0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 318 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"80E4351A76EF78185D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C4ABD86A65F13C91") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"80E4351A76EF78185D";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C4ABD86A65F13C91") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 319 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"80E4351A76EF78185D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E078DBCB76F7E408") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"80E4351A76EF78185D";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E078DBCB76F7E408") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 320 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"80E4351A76EF78185D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"955A5A28461488FC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"80E4351A76EF78185D";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"955A5A28461488FC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 321 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"80E4351A76EF78185D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E9866BE52766BDA8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"80E4351A76EF78185D";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E9866BE52766BDA8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 322 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"80E4351A76EF78185D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"57A46BABA294BCAD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"80E4351A76EF78185D";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"57A46BABA294BCAD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 323 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"80E4351A76EF78185D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C5B3F6849B5B6DFB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"80E4351A76EF78185D";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C5B3F6849B5B6DFB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 324 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"80E4351A76EF78185D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"083423D6627C12B2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"80E4351A76EF78185D";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"083423D6627C12B2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 325 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"80E4351A76EF78185D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AFA8E9E73169B29C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"80E4351A76EF78185D";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AFA8E9E73169B29C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 326 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"80E4351A76EF78185D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"458E27E50DDCC69D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"80E4351A76EF78185D";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"458E27E50DDCC69D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 327 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"80E4351A76EF78185D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1D5C45B0D21F8346") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"80E4351A76EF78185D";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1D5C45B0D21F8346") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 328 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"80E4351A76EF78185D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"079FBC2872F61A00") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"80E4351A76EF78185D";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"079FBC2872F61A00") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 329 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"80E4351A76EF78185D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1078DD4E59B3CB2E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"80E4351A76EF78185D";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1078DD4E59B3CB2E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 330 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"80E4351A76EF78185D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"12A3A637E8EDF155") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"80E4351A76EF78185D";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"000102030405060708") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"12A3A637E8EDF155") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 331 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"80E4351A76EF78185D6E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4AB3CE25A63BAE65") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"80E4351A76EF78185D6E";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4AB3CE25A63BAE65") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 332 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"80E4351A76EF78185D6E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C4CE706DC7699496") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"80E4351A76EF78185D6E";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C4CE706DC7699496") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 333 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"80E4351A76EF78185D6E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9783A25A0507F39E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"80E4351A76EF78185D6E";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9783A25A0507F39E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 334 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"80E4351A76EF78185D6E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3E57C0F611CB41BF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"80E4351A76EF78185D6E";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3E57C0F611CB41BF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 335 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"80E4351A76EF78185D6E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"80775B002B9D661C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"80E4351A76EF78185D6E";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"80775B002B9D661C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 336 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"80E4351A76EF78185D6E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2F518577E63D5867") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"80E4351A76EF78185D6E";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2F518577E63D5867") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 337 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"80E4351A76EF78185D6E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9D3388855810F677") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"80E4351A76EF78185D6E";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9D3388855810F677") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 338 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"80E4351A76EF78185D6E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F6AAE2A1340D95BA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"80E4351A76EF78185D6E";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F6AAE2A1340D95BA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 339 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"80E4351A76EF78185D6E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2C4CC0336A99D16C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"80E4351A76EF78185D6E";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2C4CC0336A99D16C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 340 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"80E4351A76EF78185D6E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8344F9B2F438C5F5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"80E4351A76EF78185D6E";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8344F9B2F438C5F5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 341 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"80E4351A76EF78185D6E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"25BDA8BADE0447DF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"80E4351A76EF78185D6E";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"25BDA8BADE0447DF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 342 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"80E4351A76EF78185D6E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9CB798A66E7FA5CB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"80E4351A76EF78185D6E";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9CB798A66E7FA5CB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 343 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"80E4351A76EF78185D6E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FCF9E43122C584B9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"80E4351A76EF78185D6E";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FCF9E43122C584B9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 344 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"80E4351A76EF78185D6E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D45602913E0E8611") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"80E4351A76EF78185D6E";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D45602913E0E8611") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 345 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"80E4351A76EF78185D6E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AF2E20A3ED26A19A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"80E4351A76EF78185D6E";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AF2E20A3ED26A19A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 346 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"80E4351A76EF78185D6E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"22A809753977D34E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"80E4351A76EF78185D6E";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"22A809753977D34E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 347 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"80E4351A76EF78185D6E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CC17AF24E7A9F69A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"80E4351A76EF78185D6E";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CC17AF24E7A9F69A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 348 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"80E4351A76EF78185D6E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EB87B752C9F63632") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"80E4351A76EF78185D6E";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EB87B752C9F63632") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 349 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"80E4351A76EF78185D6E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C7E9373720185063") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"80E4351A76EF78185D6E";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C7E9373720185063") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 350 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"80E4351A76EF78185D6E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7820DD1054B1DE21") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"80E4351A76EF78185D6E";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7820DD1054B1DE21") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 351 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"80E4351A76EF78185D6E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"95F13D6D8CF9F770") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"80E4351A76EF78185D6E";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"95F13D6D8CF9F770") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 352 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"80E4351A76EF78185D6E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B1223ECC9FFF2FE9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"80E4351A76EF78185D6E";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B1223ECC9FFF2FE9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 353 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"80E4351A76EF78185D6E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C400BF2FAF1C431D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"80E4351A76EF78185D6E";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C400BF2FAF1C431D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 354 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"80E4351A76EF78185D6E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B8DC8EE2CE6E7649") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"80E4351A76EF78185D6E";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B8DC8EE2CE6E7649") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 355 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"80E4351A76EF78185D6E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"06FE8EAC4B9C774C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"80E4351A76EF78185D6E";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"06FE8EAC4B9C774C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 356 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"80E4351A76EF78185D6E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"94E913837253A61A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"80E4351A76EF78185D6E";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"94E913837253A61A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 357 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"80E4351A76EF78185D6E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"596EC6D18B74D953") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"80E4351A76EF78185D6E";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"596EC6D18B74D953") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 358 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"80E4351A76EF78185D6E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FEF20CE0D861797D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"80E4351A76EF78185D6E";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FEF20CE0D861797D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 359 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"80E4351A76EF78185D6E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"14D4C2E2E4D40D7C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"80E4351A76EF78185D6E";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"14D4C2E2E4D40D7C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 360 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"80E4351A76EF78185D6E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4C06A0B73B1748A7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"80E4351A76EF78185D6E";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4C06A0B73B1748A7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 361 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"80E4351A76EF78185D6E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"56C5592F9BFED1E1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"80E4351A76EF78185D6E";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"56C5592F9BFED1E1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 362 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"80E4351A76EF78185D6E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"41223849B0BB00CF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"80E4351A76EF78185D6E";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"41223849B0BB00CF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 363 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"80E4351A76EF78185D6E") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"43F9433001E53AB4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"80E4351A76EF78185D6E";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"00010203040506070809") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"43F9433001E53AB4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 364 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"80E4351A76EF78185D6E1F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8A30BF994BBD98FB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"80E4351A76EF78185D6E1F";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8A30BF994BBD98FB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 365 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"80E4351A76EF78185D6E1F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"044D01D12AEFA208") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"80E4351A76EF78185D6E1F";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"044D01D12AEFA208") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 366 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"80E4351A76EF78185D6E1F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5700D3E6E881C500") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"80E4351A76EF78185D6E1F";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5700D3E6E881C500") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 367 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"80E4351A76EF78185D6E1F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FED4B14AFC4D7721") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"80E4351A76EF78185D6E1F";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FED4B14AFC4D7721") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 368 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"80E4351A76EF78185D6E1F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"40F42ABCC61B5082") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"80E4351A76EF78185D6E1F";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"40F42ABCC61B5082") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 369 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"80E4351A76EF78185D6E1F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EFD2F4CB0BBB6EF9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"80E4351A76EF78185D6E1F";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EFD2F4CB0BBB6EF9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 370 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"80E4351A76EF78185D6E1F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5DB0F939B596C0E9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"80E4351A76EF78185D6E1F";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5DB0F939B596C0E9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 371 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"80E4351A76EF78185D6E1F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3629931DD98BA324") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"80E4351A76EF78185D6E1F";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3629931DD98BA324") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 372 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"80E4351A76EF78185D6E1F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"ECCFB18F871FE7F2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"80E4351A76EF78185D6E1F";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"ECCFB18F871FE7F2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 373 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"80E4351A76EF78185D6E1F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"43C7880E19BEF36B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"80E4351A76EF78185D6E1F";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"43C7880E19BEF36B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 374 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"80E4351A76EF78185D6E1F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E53ED90633827141") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"80E4351A76EF78185D6E1F";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E53ED90633827141") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 375 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"80E4351A76EF78185D6E1F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5C34E91A83F99355") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"80E4351A76EF78185D6E1F";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5C34E91A83F99355") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 376 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"80E4351A76EF78185D6E1F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3C7A958DCF43B227") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"80E4351A76EF78185D6E1F";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3C7A958DCF43B227") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 377 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"80E4351A76EF78185D6E1F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"14D5732DD388B08F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"80E4351A76EF78185D6E1F";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"14D5732DD388B08F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 378 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"80E4351A76EF78185D6E1F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6FAD511F00A09704") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"80E4351A76EF78185D6E1F";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6FAD511F00A09704") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 379 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"80E4351A76EF78185D6E1F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E22B78C9D4F1E5D0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"80E4351A76EF78185D6E1F";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E22B78C9D4F1E5D0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 380 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"80E4351A76EF78185D6E1F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0C94DE980A2FC004") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"80E4351A76EF78185D6E1F";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0C94DE980A2FC004") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 381 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"80E4351A76EF78185D6E1F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2B04C6EE247000AC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"80E4351A76EF78185D6E1F";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2B04C6EE247000AC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 382 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"80E4351A76EF78185D6E1F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"076A468BCD9E66FD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"80E4351A76EF78185D6E1F";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"076A468BCD9E66FD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 383 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"80E4351A76EF78185D6E1F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B8A3ACACB937E8BF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"80E4351A76EF78185D6E1F";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B8A3ACACB937E8BF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 384 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"80E4351A76EF78185D6E1F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"55724CD1617FC1EE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"80E4351A76EF78185D6E1F";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"55724CD1617FC1EE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 385 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"80E4351A76EF78185D6E1F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"71A14F7072791977") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"80E4351A76EF78185D6E1F";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"71A14F7072791977") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 386 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"80E4351A76EF78185D6E1F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0483CE93429A7583") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"80E4351A76EF78185D6E1F";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0483CE93429A7583") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 387 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"80E4351A76EF78185D6E1F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"785FFF5E23E840D7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"80E4351A76EF78185D6E1F";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"785FFF5E23E840D7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 388 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"80E4351A76EF78185D6E1F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C67DFF10A61A41D2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"80E4351A76EF78185D6E1F";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C67DFF10A61A41D2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 389 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"80E4351A76EF78185D6E1F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"546A623F9FD59084") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"80E4351A76EF78185D6E1F";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"546A623F9FD59084") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 390 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"80E4351A76EF78185D6E1F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"99EDB76D66F2EFCD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"80E4351A76EF78185D6E1F";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"99EDB76D66F2EFCD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 391 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"80E4351A76EF78185D6E1F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3E717D5C35E74FE3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"80E4351A76EF78185D6E1F";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3E717D5C35E74FE3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 392 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"80E4351A76EF78185D6E1F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D457B35E09523BE2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"80E4351A76EF78185D6E1F";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D457B35E09523BE2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 393 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"80E4351A76EF78185D6E1F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8C85D10BD6917E39") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"80E4351A76EF78185D6E1F";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8C85D10BD6917E39") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 394 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"80E4351A76EF78185D6E1F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"964628937678E77F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"80E4351A76EF78185D6E1F";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"964628937678E77F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 395 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"80E4351A76EF78185D6E1F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"81A149F55D3D3651") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"80E4351A76EF78185D6E1F";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"81A149F55D3D3651") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 396 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"80E4351A76EF78185D6E1F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"837A328CEC630C2A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"80E4351A76EF78185D6E1F";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"000102030405060708090A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"837A328CEC630C2A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 397 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"80E4351A76EF78185D6E1F23") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A70929FA6BBC6DBC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"80E4351A76EF78185D6E1F23";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A70929FA6BBC6DBC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 398 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"80E4351A76EF78185D6E1F23") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"297497B20AEE574F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"80E4351A76EF78185D6E1F23";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"297497B20AEE574F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 399 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"80E4351A76EF78185D6E1F23") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7A394585C8803047") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"80E4351A76EF78185D6E1F23";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7A394585C8803047") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 400 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"80E4351A76EF78185D6E1F23") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D3ED2729DC4C8266") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"80E4351A76EF78185D6E1F23";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D3ED2729DC4C8266") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 401 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"80E4351A76EF78185D6E1F23") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6DCDBCDFE61AA5C5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"80E4351A76EF78185D6E1F23";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6DCDBCDFE61AA5C5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 402 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"80E4351A76EF78185D6E1F23") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C2EB62A82BBA9BBE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"80E4351A76EF78185D6E1F23";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C2EB62A82BBA9BBE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 403 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"80E4351A76EF78185D6E1F23") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"70896F5A959735AE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"80E4351A76EF78185D6E1F23";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"70896F5A959735AE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 404 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"80E4351A76EF78185D6E1F23") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1B10057EF98A5663") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"80E4351A76EF78185D6E1F23";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1B10057EF98A5663") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 405 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"80E4351A76EF78185D6E1F23") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C1F627ECA71E12B5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"80E4351A76EF78185D6E1F23";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C1F627ECA71E12B5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 406 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"80E4351A76EF78185D6E1F23") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6EFE1E6D39BF062C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"80E4351A76EF78185D6E1F23";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6EFE1E6D39BF062C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 407 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"80E4351A76EF78185D6E1F23") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C8074F6513838406") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"80E4351A76EF78185D6E1F23";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C8074F6513838406") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 408 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"80E4351A76EF78185D6E1F23") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"710D7F79A3F86612") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"80E4351A76EF78185D6E1F23";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"710D7F79A3F86612") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 409 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"80E4351A76EF78185D6E1F23") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"114303EEEF424760") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"80E4351A76EF78185D6E1F23";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"114303EEEF424760") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 410 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"80E4351A76EF78185D6E1F23") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"39ECE54EF38945C8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"80E4351A76EF78185D6E1F23";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"39ECE54EF38945C8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 411 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"80E4351A76EF78185D6E1F23") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4294C77C20A16243") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"80E4351A76EF78185D6E1F23";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4294C77C20A16243") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 412 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"80E4351A76EF78185D6E1F23") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CF12EEAAF4F01097") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"80E4351A76EF78185D6E1F23";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CF12EEAAF4F01097") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 413 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"80E4351A76EF78185D6E1F23") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"21AD48FB2A2E3543") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"80E4351A76EF78185D6E1F23";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"21AD48FB2A2E3543") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 414 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"80E4351A76EF78185D6E1F23") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"063D508D0471F5EB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"80E4351A76EF78185D6E1F23";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"063D508D0471F5EB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 415 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"80E4351A76EF78185D6E1F23") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2A53D0E8ED9F93BA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"80E4351A76EF78185D6E1F23";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2A53D0E8ED9F93BA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 416 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"80E4351A76EF78185D6E1F23") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"959A3ACF99361DF8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"80E4351A76EF78185D6E1F23";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"959A3ACF99361DF8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 417 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"80E4351A76EF78185D6E1F23") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"784BDAB2417E34A9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"80E4351A76EF78185D6E1F23";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"784BDAB2417E34A9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 418 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"80E4351A76EF78185D6E1F23") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5C98D9135278EC30") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"80E4351A76EF78185D6E1F23";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5C98D9135278EC30") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 419 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"80E4351A76EF78185D6E1F23") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"29BA58F0629B80C4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"80E4351A76EF78185D6E1F23";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"29BA58F0629B80C4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 420 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"80E4351A76EF78185D6E1F23") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5566693D03E9B590") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"80E4351A76EF78185D6E1F23";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5566693D03E9B590") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 421 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"80E4351A76EF78185D6E1F23") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EB446973861BB495") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"80E4351A76EF78185D6E1F23";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EB446973861BB495") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 422 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"80E4351A76EF78185D6E1F23") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7953F45CBFD465C3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"80E4351A76EF78185D6E1F23";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7953F45CBFD465C3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 423 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"80E4351A76EF78185D6E1F23") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B4D4210E46F31A8A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"80E4351A76EF78185D6E1F23";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B4D4210E46F31A8A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 424 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"80E4351A76EF78185D6E1F23") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1348EB3F15E6BAA4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"80E4351A76EF78185D6E1F23";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1348EB3F15E6BAA4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 425 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"80E4351A76EF78185D6E1F23") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F96E253D2953CEA5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"80E4351A76EF78185D6E1F23";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F96E253D2953CEA5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 426 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"80E4351A76EF78185D6E1F23") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A1BC4768F6908B7E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"80E4351A76EF78185D6E1F23";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A1BC4768F6908B7E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 427 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"80E4351A76EF78185D6E1F23") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BB7FBEF056791238") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"80E4351A76EF78185D6E1F23";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BB7FBEF056791238") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 428 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"80E4351A76EF78185D6E1F23") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AC98DF967D3CC316") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"80E4351A76EF78185D6E1F23";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AC98DF967D3CC316") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 429 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"80E4351A76EF78185D6E1F23") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AE43A4EFCC62F96D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"80E4351A76EF78185D6E1F23";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"000102030405060708090A0B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AE43A4EFCC62F96D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 430 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"80E4351A76EF78185D6E1F23BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DC661AF9F202A6E7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"80E4351A76EF78185D6E1F23BC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DC661AF9F202A6E7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 431 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"80E4351A76EF78185D6E1F23BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"521BA4B193509C14") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"80E4351A76EF78185D6E1F23BC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"521BA4B193509C14") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 432 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"80E4351A76EF78185D6E1F23BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"01567686513EFB1C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"80E4351A76EF78185D6E1F23BC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"01567686513EFB1C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 433 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"80E4351A76EF78185D6E1F23BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A882142A45F2493D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"80E4351A76EF78185D6E1F23BC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A882142A45F2493D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 434 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"80E4351A76EF78185D6E1F23BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"16A28FDC7FA46E9E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"80E4351A76EF78185D6E1F23BC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"16A28FDC7FA46E9E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 435 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"80E4351A76EF78185D6E1F23BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B98451ABB20450E5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"80E4351A76EF78185D6E1F23BC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B98451ABB20450E5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 436 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"80E4351A76EF78185D6E1F23BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0BE65C590C29FEF5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"80E4351A76EF78185D6E1F23BC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0BE65C590C29FEF5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 437 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"80E4351A76EF78185D6E1F23BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"607F367D60349D38") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"80E4351A76EF78185D6E1F23BC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"607F367D60349D38") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 438 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"80E4351A76EF78185D6E1F23BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BA9914EF3EA0D9EE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"80E4351A76EF78185D6E1F23BC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BA9914EF3EA0D9EE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 439 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"80E4351A76EF78185D6E1F23BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"15912D6EA001CD77") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"80E4351A76EF78185D6E1F23BC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"15912D6EA001CD77") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 440 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"80E4351A76EF78185D6E1F23BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B3687C668A3D4F5D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"80E4351A76EF78185D6E1F23BC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B3687C668A3D4F5D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 441 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"80E4351A76EF78185D6E1F23BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0A624C7A3A46AD49") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"80E4351A76EF78185D6E1F23BC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0A624C7A3A46AD49") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 442 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"80E4351A76EF78185D6E1F23BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6A2C30ED76FC8C3B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"80E4351A76EF78185D6E1F23BC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6A2C30ED76FC8C3B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 443 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"80E4351A76EF78185D6E1F23BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4283D64D6A378E93") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"80E4351A76EF78185D6E1F23BC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4283D64D6A378E93") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 444 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"80E4351A76EF78185D6E1F23BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"39FBF47FB91FA918") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"80E4351A76EF78185D6E1F23BC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"39FBF47FB91FA918") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 445 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"80E4351A76EF78185D6E1F23BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B47DDDA96D4EDBCC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"80E4351A76EF78185D6E1F23BC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B47DDDA96D4EDBCC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 446 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"80E4351A76EF78185D6E1F23BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5AC27BF8B390FE18") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"80E4351A76EF78185D6E1F23BC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5AC27BF8B390FE18") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 447 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"80E4351A76EF78185D6E1F23BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7D52638E9DCF3EB0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"80E4351A76EF78185D6E1F23BC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7D52638E9DCF3EB0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 448 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"80E4351A76EF78185D6E1F23BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"513CE3EB742158E1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"80E4351A76EF78185D6E1F23BC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"513CE3EB742158E1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 449 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"80E4351A76EF78185D6E1F23BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EEF509CC0088D6A3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"80E4351A76EF78185D6E1F23BC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EEF509CC0088D6A3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 450 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"80E4351A76EF78185D6E1F23BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0324E9B1D8C0FFF2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"80E4351A76EF78185D6E1F23BC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0324E9B1D8C0FFF2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 451 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"80E4351A76EF78185D6E1F23BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"27F7EA10CBC6276B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"80E4351A76EF78185D6E1F23BC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"27F7EA10CBC6276B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 452 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"80E4351A76EF78185D6E1F23BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"52D56BF3FB254B9F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"80E4351A76EF78185D6E1F23BC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"52D56BF3FB254B9F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 453 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"80E4351A76EF78185D6E1F23BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2E095A3E9A577ECB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"80E4351A76EF78185D6E1F23BC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2E095A3E9A577ECB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 454 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"80E4351A76EF78185D6E1F23BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"902B5A701FA57FCE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"80E4351A76EF78185D6E1F23BC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"902B5A701FA57FCE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 455 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"80E4351A76EF78185D6E1F23BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"023CC75F266AAE98") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"80E4351A76EF78185D6E1F23BC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"023CC75F266AAE98") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 456 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"80E4351A76EF78185D6E1F23BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CFBB120DDF4DD1D1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"80E4351A76EF78185D6E1F23BC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CFBB120DDF4DD1D1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 457 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"80E4351A76EF78185D6E1F23BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6827D83C8C5871FF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"80E4351A76EF78185D6E1F23BC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6827D83C8C5871FF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 458 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"80E4351A76EF78185D6E1F23BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8201163EB0ED05FE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"80E4351A76EF78185D6E1F23BC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8201163EB0ED05FE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 459 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"80E4351A76EF78185D6E1F23BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DAD3746B6F2E4025") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"80E4351A76EF78185D6E1F23BC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DAD3746B6F2E4025") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 460 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"80E4351A76EF78185D6E1F23BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C0108DF3CFC7D963") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"80E4351A76EF78185D6E1F23BC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C0108DF3CFC7D963") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 461 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"80E4351A76EF78185D6E1F23BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D7F7EC95E482084D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"80E4351A76EF78185D6E1F23BC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D7F7EC95E482084D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 462 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"80E4351A76EF78185D6E1F23BC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D52C97EC55DC3236") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"80E4351A76EF78185D6E1F23BC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"000102030405060708090A0B0C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D52C97EC55DC3236") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 463 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"80E4351A76EF78185D6E1F23BC42") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D3B78106CC3D730B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"80E4351A76EF78185D6E1F23BC42";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D3B78106CC3D730B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 464 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"80E4351A76EF78185D6E1F23BC42") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5DCA3F4EAD6F49F8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"80E4351A76EF78185D6E1F23BC42";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5DCA3F4EAD6F49F8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 465 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"80E4351A76EF78185D6E1F23BC42") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0E87ED796F012EF0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"80E4351A76EF78185D6E1F23BC42";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0E87ED796F012EF0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 466 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"80E4351A76EF78185D6E1F23BC42") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A7538FD57BCD9CD1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"80E4351A76EF78185D6E1F23BC42";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A7538FD57BCD9CD1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 467 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"80E4351A76EF78185D6E1F23BC42") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"19731423419BBB72") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"80E4351A76EF78185D6E1F23BC42";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"19731423419BBB72") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 468 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"80E4351A76EF78185D6E1F23BC42") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B655CA548C3B8509") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"80E4351A76EF78185D6E1F23BC42";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B655CA548C3B8509") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 469 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"80E4351A76EF78185D6E1F23BC42") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0437C7A632162B19") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"80E4351A76EF78185D6E1F23BC42";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0437C7A632162B19") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 470 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"80E4351A76EF78185D6E1F23BC42") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6FAEAD825E0B48D4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"80E4351A76EF78185D6E1F23BC42";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6FAEAD825E0B48D4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 471 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"80E4351A76EF78185D6E1F23BC42") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B5488F10009F0C02") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"80E4351A76EF78185D6E1F23BC42";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B5488F10009F0C02") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 472 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"80E4351A76EF78185D6E1F23BC42") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1A40B6919E3E189B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"80E4351A76EF78185D6E1F23BC42";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1A40B6919E3E189B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 473 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"80E4351A76EF78185D6E1F23BC42") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BCB9E799B4029AB1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"80E4351A76EF78185D6E1F23BC42";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BCB9E799B4029AB1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 474 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"80E4351A76EF78185D6E1F23BC42") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"05B3D785047978A5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"80E4351A76EF78185D6E1F23BC42";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"05B3D785047978A5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 475 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"80E4351A76EF78185D6E1F23BC42") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"65FDAB1248C359D7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"80E4351A76EF78185D6E1F23BC42";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"65FDAB1248C359D7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 476 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"80E4351A76EF78185D6E1F23BC42") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4D524DB254085B7F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"80E4351A76EF78185D6E1F23BC42";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4D524DB254085B7F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 477 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"80E4351A76EF78185D6E1F23BC42") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"362A6F8087207CF4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"80E4351A76EF78185D6E1F23BC42";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"362A6F8087207CF4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 478 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"80E4351A76EF78185D6E1F23BC42") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BBAC465653710E20") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"80E4351A76EF78185D6E1F23BC42";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BBAC465653710E20") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 479 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"80E4351A76EF78185D6E1F23BC42") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5513E0078DAF2BF4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"80E4351A76EF78185D6E1F23BC42";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5513E0078DAF2BF4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 480 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"80E4351A76EF78185D6E1F23BC42") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7283F871A3F0EB5C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"80E4351A76EF78185D6E1F23BC42";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7283F871A3F0EB5C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 481 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"80E4351A76EF78185D6E1F23BC42") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5EED78144A1E8D0D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"80E4351A76EF78185D6E1F23BC42";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5EED78144A1E8D0D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 482 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"80E4351A76EF78185D6E1F23BC42") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E12492333EB7034F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"80E4351A76EF78185D6E1F23BC42";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E12492333EB7034F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 483 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"80E4351A76EF78185D6E1F23BC42") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0CF5724EE6FF2A1E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"80E4351A76EF78185D6E1F23BC42";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0CF5724EE6FF2A1E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 484 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"80E4351A76EF78185D6E1F23BC42") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"282671EFF5F9F287") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"80E4351A76EF78185D6E1F23BC42";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"282671EFF5F9F287") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 485 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"80E4351A76EF78185D6E1F23BC42") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5D04F00CC51A9E73") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"80E4351A76EF78185D6E1F23BC42";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5D04F00CC51A9E73") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 486 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"80E4351A76EF78185D6E1F23BC42") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"21D8C1C1A468AB27") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"80E4351A76EF78185D6E1F23BC42";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"21D8C1C1A468AB27") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 487 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"80E4351A76EF78185D6E1F23BC42") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9FFAC18F219AAA22") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"80E4351A76EF78185D6E1F23BC42";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9FFAC18F219AAA22") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 488 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"80E4351A76EF78185D6E1F23BC42") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0DED5CA018557B74") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"80E4351A76EF78185D6E1F23BC42";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0DED5CA018557B74") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 489 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"80E4351A76EF78185D6E1F23BC42") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C06A89F2E172043D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"80E4351A76EF78185D6E1F23BC42";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C06A89F2E172043D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 490 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"80E4351A76EF78185D6E1F23BC42") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"67F643C3B267A413") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"80E4351A76EF78185D6E1F23BC42";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"67F643C3B267A413") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 491 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"80E4351A76EF78185D6E1F23BC42") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8DD08DC18ED2D012") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"80E4351A76EF78185D6E1F23BC42";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8DD08DC18ED2D012") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 492 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"80E4351A76EF78185D6E1F23BC42") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D502EF94511195C9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"80E4351A76EF78185D6E1F23BC42";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D502EF94511195C9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 493 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"80E4351A76EF78185D6E1F23BC42") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CFC1160CF1F80C8F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"80E4351A76EF78185D6E1F23BC42";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CFC1160CF1F80C8F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 494 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"80E4351A76EF78185D6E1F23BC42") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D826776ADABDDDA1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"80E4351A76EF78185D6E1F23BC42";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D826776ADABDDDA1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 495 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"80E4351A76EF78185D6E1F23BC42") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DAFD0C136BE3E7DA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"80E4351A76EF78185D6E1F23BC42";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"000102030405060708090A0B0C0D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DAFD0C136BE3E7DA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 496 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"80E4351A76EF78185D6E1F23BC42D0") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"777DE81E009C1430") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"80E4351A76EF78185D6E1F23BC42D0";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"777DE81E009C1430") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 497 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"80E4351A76EF78185D6E1F23BC42D0") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F900565661CE2EC3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"80E4351A76EF78185D6E1F23BC42D0";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F900565661CE2EC3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 498 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"80E4351A76EF78185D6E1F23BC42D0") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AA4D8461A3A049CB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"80E4351A76EF78185D6E1F23BC42D0";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AA4D8461A3A049CB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 499 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"80E4351A76EF78185D6E1F23BC42D0") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0399E6CDB76CFBEA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B0C0D0E0F";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"80E4351A76EF78185D6E1F23BC42D0";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0399E6CDB76CFBEA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --======================================================================================= 

      wait;
   end process;

END;
