--
-- SKINNY-AEAD Reference Hardware Implementation
-- 
-- Copyright 2019:
--     Amir Moradi & Pascal Sasdrich for the SKINNY Team
--     https://sites.google.com/site/skinnycipher/
-- 
-- This program is free software; you can redistribute it and/or
-- modify it under the terms of the GNU General Public License as
-- published by the Free Software Foundation; either version 2 of the
-- License, or (at your option) any later version.
-- 
-- This program is distributed in the hope that it will be useful, but
-- WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE. See the GNU
-- General Public License for more details.
-- 

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
ENTITY SKINNY_tk2_AEAD_M5_Test_Part2 IS
END SKINNY_tk2_AEAD_M5_Test_Part2;
 
ARCHITECTURE behavior OF SKINNY_tk2_AEAD_M5_Test_Part2 IS 
 
	constant tl		 : integer := 0; -- 128-bit tag -> M5
 
 
   COMPONENT SKINNY_tk2_AEAD
	Generic (
		tl				 : integer); -- 0: 128-bit tag,   1: 64-bit tag
	Port (  
		clk          : in  STD_LOGIC;
		rst      	 : in  STD_LOGIC;
		a_data       : in  STD_LOGIC;
		enc          : in  STD_LOGIC;
		dec          : in  STD_LOGIC;
		gen_tag      : in  std_logic;
		Input        : in  STD_LOGIC_VECTOR (127 downto 0);  -- Message or Associated Data
		N            : in  STD_LOGIC_VECTOR ( 95 downto 0);
		K            : in  STD_LOGIC_VECTOR (127 downto 0);
		Block_Size	 : in  STD_LOGIC_VECTOR (  3 downto 0); -- Size of the given block as Input (in BYTES) - 1
		Output       : out STD_LOGIC_VECTOR (127 downto 0); -- Ciphertext or Plaintext
		Tag			 : out STD_LOGIC_VECTOR (127-tl*64 downto 0); -- Tag
		done         : out STD_LOGIC);
   END COMPONENT;
    

   --Inputs
   signal clk 			: std_logic := '0';
   signal rst 			: std_logic := '0';
   signal a_data 		: std_logic := '0';
   signal enc 			: std_logic := '0';
   signal dec 			: std_logic := '0';
   signal gen_tag 	: std_logic := '0';
   signal Input 		: std_logic_vector(127 downto 0) := (others => '0');
   signal N 			: std_logic_vector( 95 downto 0) := (others => '0');
   signal K 			: std_logic_vector(127 downto 0) := (others => '0');
   signal Block_Size : std_logic_vector(  3 downto 0) := (others => '0');

 	--Outputs
   signal Output 		: std_logic_vector(127 downto 0);
   signal Tag 		   : std_logic_vector(127-tl*64 downto 0);
   signal done 		: std_logic;

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
   uut: SKINNY_tk2_AEAD 
	GENERIC MAP (
		tl => tl)
	PORT MAP (
		clk 			=> clk,
		rst 			=> rst,
		a_data 		=> a_data,
		enc 			=> enc,
		dec 			=> dec,
		gen_tag 		=> gen_tag,
		Input 		=> Input,
		N 				=> N,
		K 				=> K,
		Block_Size 	=> Block_Size,
		Output 		=> Output,
		Tag			=> Tag,
		done 			=> done
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      --------- test no. 500 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"684E406EF1682AE8A1E5093C8539C0") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"52836243399834AA06ACDC1AF68533E9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"684E406EF1682AE8A1E5093C8539C0";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"52836243399834AA06ACDC1AF68533E9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 501 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"684E406EF1682AE8A1E5093C8539C0") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"703119B1449D130F50AA31110FA25506") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"684E406EF1682AE8A1E5093C8539C0";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"703119B1449D130F50AA31110FA25506") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 502 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"684E406EF1682AE8A1E5093C8539C0") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E540E45F9981DDAEF6B958533053C745") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"684E406EF1682AE8A1E5093C8539C0";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E540E45F9981DDAEF6B958533053C745") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 503 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"684E406EF1682AE8A1E5093C8539C0") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"54D0E8475FCEEC15A94AA77EDAF4485D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"684E406EF1682AE8A1E5093C8539C0";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"54D0E8475FCEEC15A94AA77EDAF4485D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 504 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"684E406EF1682AE8A1E5093C8539C0") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E7D828AB368AF3F46EACCB77CE3BE28F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"684E406EF1682AE8A1E5093C8539C0";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E7D828AB368AF3F46EACCB77CE3BE28F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 505 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"684E406EF1682AE8A1E5093C8539C0") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3BD443232E95B2A30A5B5C7B6CDC1216") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"684E406EF1682AE8A1E5093C8539C0";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3BD443232E95B2A30A5B5C7B6CDC1216") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 506 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"684E406EF1682AE8A1E5093C8539C0") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8BCC9879F832BBE24B619B79F330882D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"684E406EF1682AE8A1E5093C8539C0";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8BCC9879F832BBE24B619B79F330882D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 507 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"684E406EF1682AE8A1E5093C8539C0") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F4C3712D047044C1C0F4F7F19243A349") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"684E406EF1682AE8A1E5093C8539C0";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F4C3712D047044C1C0F4F7F19243A349") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 508 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"684E406EF1682AE8A1E5093C8539C0") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6F06B992E63A6B14B2EE650A10DDE8EB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"684E406EF1682AE8A1E5093C8539C0";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6F06B992E63A6B14B2EE650A10DDE8EB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 509 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"684E406EF1682AE8A1E5093C8539C0") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"03BE39A6518CFBFAC2DEC5A604F5810E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"684E406EF1682AE8A1E5093C8539C0";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"03BE39A6518CFBFAC2DEC5A604F5810E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 510 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"684E406EF1682AE8A1E5093C8539C0") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5CDA94DF4CA880CDE7B2AEE6A39DF6CB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"684E406EF1682AE8A1E5093C8539C0";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5CDA94DF4CA880CDE7B2AEE6A39DF6CB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 511 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"684E406EF1682AE8A1E5093C8539C0") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1A9EE7DD508A2A087D12994ACDBF723D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"684E406EF1682AE8A1E5093C8539C0";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1A9EE7DD508A2A087D12994ACDBF723D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 512 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"684E406EF1682AE8A1E5093C8539C0") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BFB8DB2499CAB9DC764757292B9C43B9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"684E406EF1682AE8A1E5093C8539C0";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BFB8DB2499CAB9DC764757292B9C43B9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 513 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"684E406EF1682AE8A1E5093C8539C0") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A5C93A2343410E098C3A1603A0A5BC85") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"684E406EF1682AE8A1E5093C8539C0";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A5C93A2343410E098C3A1603A0A5BC85") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 514 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"684E406EF1682AE8A1E5093C8539C0") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D428A794DA78A23AF4C123065302CB04") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"684E406EF1682AE8A1E5093C8539C0";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D428A794DA78A23AF4C123065302CB04") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 515 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"684E406EF1682AE8A1E5093C8539C0") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1E652B8A72D3D4D1847500425227BA71") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"684E406EF1682AE8A1E5093C8539C0";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1E652B8A72D3D4D1847500425227BA71") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 516 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"684E406EF1682AE8A1E5093C8539C0") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"96E4D1D98BE9D6521C26F48C89D36520") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"684E406EF1682AE8A1E5093C8539C0";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"96E4D1D98BE9D6521C26F48C89D36520") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 517 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"684E406EF1682AE8A1E5093C8539C0") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8ABAB1C16D143D05C35CE7EE824AD3D3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"684E406EF1682AE8A1E5093C8539C0";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8ABAB1C16D143D05C35CE7EE824AD3D3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 518 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"684E406EF1682AE8A1E5093C8539C0") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7B6C837D6B7EA6DC59E0CF510F5BD228") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"684E406EF1682AE8A1E5093C8539C0";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7B6C837D6B7EA6DC59E0CF510F5BD228") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 519 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"684E406EF1682AE8A1E5093C8539C0") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7412A4008002483D1AF85EE573A5510D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"684E406EF1682AE8A1E5093C8539C0";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7412A4008002483D1AF85EE573A5510D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 520 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"684E406EF1682AE8A1E5093C8539C0") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"92B9157C19A26BD4CA7C9A84B53CD303") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"684E406EF1682AE8A1E5093C8539C0";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"92B9157C19A26BD4CA7C9A84B53CD303") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 521 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"684E406EF1682AE8A1E5093C8539C0") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"501B26BF8568244C426D04EF82E69833") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"684E406EF1682AE8A1E5093C8539C0";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"501B26BF8568244C426D04EF82E69833") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 522 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"684E406EF1682AE8A1E5093C8539C0") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F4D7F6917F8C82B5E471A09B5624AAB0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"684E406EF1682AE8A1E5093C8539C0";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F4D7F6917F8C82B5E471A09B5624AAB0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 523 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"684E406EF1682AE8A1E5093C8539C0") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"16B8C48CA4CD71B5EEFE4CE8D43993E6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"684E406EF1682AE8A1E5093C8539C0";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"16B8C48CA4CD71B5EEFE4CE8D43993E6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 524 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"684E406EF1682AE8A1E5093C8539C0") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6A9E9D9A8406918CC06F2934F0C5A8D2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"684E406EF1682AE8A1E5093C8539C0";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6A9E9D9A8406918CC06F2934F0C5A8D2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 525 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"684E406EF1682AE8A1E5093C8539C0") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7D19D87C0F88525424358DA2C709693C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"684E406EF1682AE8A1E5093C8539C0";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7D19D87C0F88525424358DA2C709693C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 526 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"684E406EF1682AE8A1E5093C8539C0") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"853713269B01FA0C477B004152E2D9AE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"684E406EF1682AE8A1E5093C8539C0";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"853713269B01FA0C477B004152E2D9AE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 527 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"684E406EF1682AE8A1E5093C8539C0") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D1039E43B5CA36BF113A305A554990C2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"684E406EF1682AE8A1E5093C8539C0";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D1039E43B5CA36BF113A305A554990C2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 528 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"684E406EF1682AE8A1E5093C8539C0") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"376E24FDC1A34B1FE6F40359F016754F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"684E406EF1682AE8A1E5093C8539C0";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"000102030405060708090A0B0C0D0E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"376E24FDC1A34B1FE6F40359F016754F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 529 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0E49D046AE510C840C9B74289FBBB533") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0E49D046AE510C840C9B74289FBBB533") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 530 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F8C55013CA4ED4CBEB91FEF049FC6610") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F8C55013CA4ED4CBEB91FEF049FC6610") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 531 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7580DD8480FA9149963B9FE5C5EC4112") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7580DD8480FA9149963B9FE5C5EC4112") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 532 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A16DE968DBEB3BF2373D659EE1F7F183") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A16DE968DBEB3BF2373D659EE1F7F183") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 533 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3020F15212773AFFD0985DDE70803D6C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3020F15212773AFFD0985DDE70803D6C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 534 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"12928AA06F721D5A869EB0D589A75B83") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"12928AA06F721D5A869EB0D589A75B83") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 535 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"87E3774EB26ED3FB208DD997B656C9C0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"87E3774EB26ED3FB208DD997B656C9C0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 536 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"36737B567421E2407F7E26BA5CF146D8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"36737B567421E2407F7E26BA5CF146D8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 537 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"857BBBBA1D65FDA1B8984AB3483EEC0A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"857BBBBA1D65FDA1B8984AB3483EEC0A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 538 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5977D032057ABCF6DC6FDDBFEAD91C93") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5977D032057ABCF6DC6FDDBFEAD91C93") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 539 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E96F0B68D3DDB5B79D551ABD753586A8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E96F0B68D3DDB5B79D551ABD753586A8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 540 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9660E23C2F9F4A9416C076351446ADCC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9660E23C2F9F4A9416C076351446ADCC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 541 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0DA52A83CDD5654164DAE4CE96D8E66E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0DA52A83CDD5654164DAE4CE96D8E66E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 542 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"611DAAB77A63F5AF14EA446282F08F8B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"611DAAB77A63F5AF14EA446282F08F8B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 543 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3E7907CE67478E9831862F222598F84E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3E7907CE67478E9831862F222598F84E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 544 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"783D74CC7B65245DAB26188E4BBA7CB8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"783D74CC7B65245DAB26188E4BBA7CB8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 545 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DD1B4835B225B789A073D6EDAD994D3C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DD1B4835B225B789A073D6EDAD994D3C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 546 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C76AA93268AE005C5A0E97C726A0B200") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C76AA93268AE005C5A0E97C726A0B200") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 547 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B68B3485F197AC6F22F5A2C2D507C581") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B68B3485F197AC6F22F5A2C2D507C581") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 548 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7CC6B89B593CDA8452418186D422B4F4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7CC6B89B593CDA8452418186D422B4F4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 549 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F44742C8A006D807CA1275480FD66BA5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F44742C8A006D807CA1275480FD66BA5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 550 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E81922D046FB33501568662A044FDD56") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E81922D046FB33501568662A044FDD56") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 551 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"19CF106C4091A8898FD44E95895EDCAD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"19CF106C4091A8898FD44E95895EDCAD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 552 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"16B13711ABED4668CCCCDF21F5A05F88") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"16B13711ABED4668CCCCDF21F5A05F88") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 553 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F01A866D324D65811C481B403339DD86") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F01A866D324D65811C481B403339DD86") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 554 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"32B8B5AEAE872A199459852B04E396B6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"32B8B5AEAE872A199459852B04E396B6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 555 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9674658054638CE03245215FD021A435") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9674658054638CE03245215FD021A435") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 556 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"741B579D8F227FE038CACD2C523C9D63") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"741B579D8F227FE038CACD2C523C9D63") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 557 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"083D0E8BAFE99FD9165BA8F076C0A657") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"083D0E8BAFE99FD9165BA8F076C0A657") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 558 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1FBA4B6D24675C01F2010C66410C67B9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1FBA4B6D24675C01F2010C66410C67B9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 559 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E7948037B0EEF459914F8185D4E7D72B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E7948037B0EEF459914F8185D4E7D72B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 560 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B3A00D529E2538EAC70EB19ED34C9E47") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B3A00D529E2538EAC70EB19ED34C9E47") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 561 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"55CDB7ECEA4C454A30C0829D76137BCA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"55CDB7ECEA4C454A30C0829D76137BCA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 562 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"46") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0A0F4CF8346DF50C55C1C50837C9A8AF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"46";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0A0F4CF8346DF50C55C1C50837C9A8AF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 563 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"46") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FC83CCAD50722D43B2CB4FD0E18E7B8C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"46";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FC83CCAD50722D43B2CB4FD0E18E7B8C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 564 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"46") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"71C6413A1AC668C1CF612EC56D9E5C8E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"46";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"71C6413A1AC668C1CF612EC56D9E5C8E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 565 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"46") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A52B75D641D7C27A6E67D4BE4985EC1F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"46";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A52B75D641D7C27A6E67D4BE4985EC1F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 566 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"46") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"34666DEC884BC37789C2ECFED8F220F0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"46";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"34666DEC884BC37789C2ECFED8F220F0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 567 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"46") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"16D4161EF54EE4D2DFC401F521D5461F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"46";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"16D4161EF54EE4D2DFC401F521D5461F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 568 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"46") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"83A5EBF028522A7379D768B71E24D45C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"46";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"83A5EBF028522A7379D768B71E24D45C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 569 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"46") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3235E7E8EE1D1BC82624979AF4835B44") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"46";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3235E7E8EE1D1BC82624979AF4835B44") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 570 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"46") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"813D270487590429E1C2FB93E04CF196") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"46";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"813D270487590429E1C2FB93E04CF196") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 571 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"46") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5D314C8C9F46457E85356C9F42AB010F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"46";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5D314C8C9F46457E85356C9F42AB010F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 572 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"46") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"ED2997D649E14C3FC40FAB9DDD479B34") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"46";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"ED2997D649E14C3FC40FAB9DDD479B34") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 573 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"46") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"92267E82B5A3B31C4F9AC715BC34B050") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"46";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"92267E82B5A3B31C4F9AC715BC34B050") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 574 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"46") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"09E3B63D57E99CC93D8055EE3EAAFBF2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"46";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"09E3B63D57E99CC93D8055EE3EAAFBF2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 575 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"46") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"655B3609E05F0C274DB0F5422A829217") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"46";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"655B3609E05F0C274DB0F5422A829217") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 576 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"46") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3A3F9B70FD7B771068DC9E028DEAE5D2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"46";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3A3F9B70FD7B771068DC9E028DEAE5D2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 577 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"46") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7C7BE872E159DDD5F27CA9AEE3C86124") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"46";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7C7BE872E159DDD5F27CA9AEE3C86124") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 578 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"46") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D95DD48B28194E01F92967CD05EB50A0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"46";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D95DD48B28194E01F92967CD05EB50A0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 579 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"46") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C32C358CF292F9D4035426E78ED2AF9C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"46";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C32C358CF292F9D4035426E78ED2AF9C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 580 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"46") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B2CDA83B6BAB55E77BAF13E27D75D81D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"46";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B2CDA83B6BAB55E77BAF13E27D75D81D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 581 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"46") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"78802425C300230C0B1B30A67C50A968") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"46";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"78802425C300230C0B1B30A67C50A968") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 582 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"46") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F001DE763A3A218F9348C468A7A47639") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"46";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F001DE763A3A218F9348C468A7A47639") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 583 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"46") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EC5FBE6EDCC7CAD84C32D70AAC3DC0CA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"46";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EC5FBE6EDCC7CAD84C32D70AAC3DC0CA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 584 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"46") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1D898CD2DAAD5101D68EFFB5212CC131") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"46";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1D898CD2DAAD5101D68EFFB5212CC131") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 585 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"46") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"12F7ABAF31D1BFE095966E015DD24214") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"46";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"12F7ABAF31D1BFE095966E015DD24214") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 586 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"46") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F45C1AD3A8719C094512AA609B4BC01A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"46";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F45C1AD3A8719C094512AA609B4BC01A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 587 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"46") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"36FE291034BBD391CD03340BAC918B2A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"46";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"36FE291034BBD391CD03340BAC918B2A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 588 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"46") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9232F93ECE5F75686B1F907F7853B9A9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"46";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9232F93ECE5F75686B1F907F7853B9A9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 589 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"46") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"705DCB23151E866861907C0CFA4E80FF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"46";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"705DCB23151E866861907C0CFA4E80FF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 590 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"46") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0C7B923535D566514F0119D0DEB2BBCB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"46";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0C7B923535D566514F0119D0DEB2BBCB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 591 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"46") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1BFCD7D3BE5BA589AB5BBD46E97E7A25") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"46";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1BFCD7D3BE5BA589AB5BBD46E97E7A25") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 592 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"46") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E3D21C892AD20DD1C81530A57C95CAB7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"46";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E3D21C892AD20DD1C81530A57C95CAB7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 593 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"46") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B7E691EC0419C1629E5400BE7B3E83DB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"46";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B7E691EC0419C1629E5400BE7B3E83DB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 594 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"46") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"518B2B527070BCC2699A33BDDE616656") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"46";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-0)) = x"10") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"518B2B527070BCC2699A33BDDE616656") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 595 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"46AB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C160D3E3F09D185A61C351A48DEDE877") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"46AB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C160D3E3F09D185A61C351A48DEDE877") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 596 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"46AB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"37EC53B69482C01586C9DB7C5BAA3B54") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"46AB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"37EC53B69482C01586C9DB7C5BAA3B54") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 597 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"46AB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BAA9DE21DE368597FB63BA69D7BA1C56") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"46AB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BAA9DE21DE368597FB63BA69D7BA1C56") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 598 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"46AB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6E44EACD85272F2C5A654012F3A1ACC7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"46AB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6E44EACD85272F2C5A654012F3A1ACC7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 599 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"46AB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FF09F2F74CBB2E21BDC0785262D66028") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"46AB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FF09F2F74CBB2E21BDC0785262D66028") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 600 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"46AB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DDBB890531BE0984EBC695599BF106C7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"46AB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DDBB890531BE0984EBC695599BF106C7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 601 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"46AB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"48CA74EBECA2C7254DD5FC1BA4009484") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"46AB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"48CA74EBECA2C7254DD5FC1BA4009484") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 602 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"46AB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F95A78F32AEDF69E122603364EA71B9C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"46AB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F95A78F32AEDF69E122603364EA71B9C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 603 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"46AB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4A52B81F43A9E97FD5C06F3F5A68B14E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"46AB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4A52B81F43A9E97FD5C06F3F5A68B14E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 604 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"46AB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"965ED3975BB6A828B137F833F88F41D7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"46AB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"965ED3975BB6A828B137F833F88F41D7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 605 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"46AB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"264608CD8D11A169F00D3F316763DBEC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"46AB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"264608CD8D11A169F00D3F316763DBEC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 606 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"46AB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5949E19971535E4A7B9853B90610F088") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"46AB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5949E19971535E4A7B9853B90610F088") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 607 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"46AB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C28C29269319719F0982C142848EBB2A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"46AB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C28C29269319719F0982C142848EBB2A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 608 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"46AB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AE34A91224AFE17179B261EE90A6D2CF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"46AB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AE34A91224AFE17179B261EE90A6D2CF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 609 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"46AB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F150046B398B9A465CDE0AAE37CEA50A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"46AB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F150046B398B9A465CDE0AAE37CEA50A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 610 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"46AB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B714776925A93083C67E3D0259EC21FC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"46AB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B714776925A93083C67E3D0259EC21FC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 611 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"46AB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"12324B90ECE9A357CD2BF361BFCF1078") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"46AB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"12324B90ECE9A357CD2BF361BFCF1078") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 612 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"46AB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0843AA97366214823756B24B34F6EF44") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"46AB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0843AA97366214823756B24B34F6EF44") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 613 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"46AB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"79A23720AF5BB8B14FAD874EC75198C5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"46AB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"79A23720AF5BB8B14FAD874EC75198C5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 614 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"46AB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B3EFBB3E07F0CE5A3F19A40AC674E9B0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"46AB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B3EFBB3E07F0CE5A3F19A40AC674E9B0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 615 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"46AB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3B6E416DFECACCD9A74A50C41D8036E1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"46AB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3B6E416DFECACCD9A74A50C41D8036E1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 616 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"46AB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"273021751837278E783043A616198012") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"46AB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"273021751837278E783043A616198012") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 617 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"46AB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D6E613C91E5DBC57E28C6B199B0881E9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"46AB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D6E613C91E5DBC57E28C6B199B0881E9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 618 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"46AB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D99834B4F52152B6A194FAADE7F602CC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"46AB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D99834B4F52152B6A194FAADE7F602CC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 619 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"46AB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3F3385C86C81715F71103ECC216F80C2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"46AB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3F3385C86C81715F71103ECC216F80C2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 620 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"46AB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FD91B60BF04B3EC7F901A0A716B5CBF2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"46AB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FD91B60BF04B3EC7F901A0A716B5CBF2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 621 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"46AB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"595D66250AAF983E5F1D04D3C277F971") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"46AB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"595D66250AAF983E5F1D04D3C277F971") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 622 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"46AB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BB325438D1EE6B3E5592E8A0406AC027") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"46AB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BB325438D1EE6B3E5592E8A0406AC027") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 623 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"46AB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C7140D2EF1258B077B038D7C6496FB13") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"46AB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C7140D2EF1258B077B038D7C6496FB13") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 624 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"46AB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D09348C87AAB48DF9F5929EA535A3AFD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"46AB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D09348C87AAB48DF9F5929EA535A3AFD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 625 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"46AB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"28BD8392EE22E087FC17A409C6B18A6F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"46AB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"28BD8392EE22E087FC17A409C6B18A6F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 626 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"46AB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7C890EF7C0E92C34AA569412C11AC303") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"46AB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7C890EF7C0E92C34AA569412C11AC303") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 627 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"46AB") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9AE4B449B48051945D98A7116445268E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"46AB";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-1)) = x"1011") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9AE4B449B48051945D98A7116445268E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 628 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"46AB5D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"12F85BF5D2E0EA46BC8BFAE644BEB841") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"46AB5D";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"12F85BF5D2E0EA46BC8BFAE644BEB841") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 629 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"46AB5D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E474DBA0B6FF32095B81703E92F96B62") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"46AB5D";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E474DBA0B6FF32095B81703E92F96B62") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 630 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"46AB5D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"69315637FC4B778B262B112B1EE94C60") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"46AB5D";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"69315637FC4B778B262B112B1EE94C60") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 631 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"46AB5D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BDDC62DBA75ADD30872DEB503AF2FCF1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"46AB5D";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BDDC62DBA75ADD30872DEB503AF2FCF1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 632 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"46AB5D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2C917AE16EC6DC3D6088D310AB85301E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"46AB5D";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2C917AE16EC6DC3D6088D310AB85301E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 633 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"46AB5D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0E23011313C3FB98368E3E1B52A256F1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"46AB5D";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0E23011313C3FB98368E3E1B52A256F1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 634 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"46AB5D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9B52FCFDCEDF3539909D57596D53C4B2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"46AB5D";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9B52FCFDCEDF3539909D57596D53C4B2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 635 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"46AB5D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2AC2F0E508900482CF6EA87487F44BAA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"46AB5D";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2AC2F0E508900482CF6EA87487F44BAA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 636 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"46AB5D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"99CA300961D41B630888C47D933BE178") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"46AB5D";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"99CA300961D41B630888C47D933BE178") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 637 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"46AB5D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"45C65B8179CB5A346C7F537131DC11E1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"46AB5D";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"45C65B8179CB5A346C7F537131DC11E1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 638 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"46AB5D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F5DE80DBAF6C53752D459473AE308BDA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"46AB5D";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F5DE80DBAF6C53752D459473AE308BDA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 639 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"46AB5D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8AD1698F532EAC56A6D0F8FBCF43A0BE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"46AB5D";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8AD1698F532EAC56A6D0F8FBCF43A0BE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 640 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"46AB5D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1114A130B1648383D4CA6A004DDDEB1C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"46AB5D";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1114A130B1648383D4CA6A004DDDEB1C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 641 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"46AB5D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7DAC210406D2136DA4FACAAC59F582F9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"46AB5D";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7DAC210406D2136DA4FACAAC59F582F9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 642 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"46AB5D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"22C88C7D1BF6685A8196A1ECFE9DF53C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"46AB5D";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"22C88C7D1BF6685A8196A1ECFE9DF53C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 643 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"46AB5D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"648CFF7F07D4C29F1B36964090BF71CA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"46AB5D";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"648CFF7F07D4C29F1B36964090BF71CA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 644 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"46AB5D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C1AAC386CE94514B10635823769C404E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"46AB5D";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C1AAC386CE94514B10635823769C404E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 645 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"46AB5D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DBDB2281141FE69EEA1E1909FDA5BF72") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"46AB5D";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DBDB2281141FE69EEA1E1909FDA5BF72") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 646 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"46AB5D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AA3ABF368D264AAD92E52C0C0E02C8F3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"46AB5D";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AA3ABF368D264AAD92E52C0C0E02C8F3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 647 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"46AB5D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"60773328258D3C46E2510F480F27B986") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"46AB5D";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"60773328258D3C46E2510F480F27B986") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 648 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"46AB5D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E8F6C97BDCB73EC57A02FB86D4D366D7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"46AB5D";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E8F6C97BDCB73EC57A02FB86D4D366D7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 649 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"46AB5D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F4A8A9633A4AD592A578E8E4DF4AD024") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"46AB5D";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F4A8A9633A4AD592A578E8E4DF4AD024") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 650 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"46AB5D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"057E9BDF3C204E4B3FC4C05B525BD1DF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"46AB5D";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"057E9BDF3C204E4B3FC4C05B525BD1DF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 651 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"46AB5D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0A00BCA2D75CA0AA7CDC51EF2EA552FA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"46AB5D";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0A00BCA2D75CA0AA7CDC51EF2EA552FA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 652 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"46AB5D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"ECAB0DDE4EFC8343AC58958EE83CD0F4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"46AB5D";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"ECAB0DDE4EFC8343AC58958EE83CD0F4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 653 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"46AB5D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2E093E1DD236CCDB24490BE5DFE69BC4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"46AB5D";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2E093E1DD236CCDB24490BE5DFE69BC4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 654 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"46AB5D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8AC5EE3328D26A228255AF910B24A947") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"46AB5D";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8AC5EE3328D26A228255AF910B24A947") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 655 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"46AB5D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"68AADC2EF393992288DA43E289399011") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"46AB5D";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"68AADC2EF393992288DA43E289399011") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 656 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"46AB5D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"148C8538D358791BA64B263EADC5AB25") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"46AB5D";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"148C8538D358791BA64B263EADC5AB25") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 657 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"46AB5D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"030BC0DE58D6BAC3421182A89A096ACB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"46AB5D";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"030BC0DE58D6BAC3421182A89A096ACB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 658 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"46AB5D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FB250B84CC5F129B215F0F4B0FE2DA59") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"46AB5D";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FB250B84CC5F129B215F0F4B0FE2DA59") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 659 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"46AB5D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AF1186E1E294DE28771E3F5008499335") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"46AB5D";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AF1186E1E294DE28771E3F5008499335") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 660 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"46AB5D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"497C3C5F96FDA38880D00C53AD1676B8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"46AB5D";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-2)) = x"101112") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"497C3C5F96FDA38880D00C53AD1676B8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 661 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"46AB5D56") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BFDFF01136FE0F62A607599FD1312F8E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"46AB5D56";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BFDFF01136FE0F62A607599FD1312F8E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 662 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"46AB5D56") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4953704452E1D72D410DD3470776FCAD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"46AB5D56";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4953704452E1D72D410DD3470776FCAD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 663 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"46AB5D56") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C416FDD3185592AF3CA7B2528B66DBAF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"46AB5D56";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C416FDD3185592AF3CA7B2528B66DBAF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 664 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"46AB5D56") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"10FBC93F434438149DA14829AF7D6B3E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"46AB5D56";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"10FBC93F434438149DA14829AF7D6B3E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 665 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"46AB5D56") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"81B6D1058AD839197A0470693E0AA7D1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"46AB5D56";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"81B6D1058AD839197A0470693E0AA7D1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 666 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"46AB5D56") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A304AAF7F7DD1EBC2C029D62C72DC13E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"46AB5D56";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A304AAF7F7DD1EBC2C029D62C72DC13E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 667 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"46AB5D56") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"367557192AC1D01D8A11F420F8DC537D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"46AB5D56";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"367557192AC1D01D8A11F420F8DC537D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 668 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"46AB5D56") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"87E55B01EC8EE1A6D5E20B0D127BDC65") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"46AB5D56";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"87E55B01EC8EE1A6D5E20B0D127BDC65") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 669 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"46AB5D56") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"34ED9BED85CAFE471204670406B476B7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"46AB5D56";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"34ED9BED85CAFE471204670406B476B7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 670 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"46AB5D56") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E8E1F0659DD5BF1076F3F008A453862E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"46AB5D56";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E8E1F0659DD5BF1076F3F008A453862E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 671 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"46AB5D56") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"58F92B3F4B72B65137C9370A3BBF1C15") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"46AB5D56";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"58F92B3F4B72B65137C9370A3BBF1C15") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 672 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"46AB5D56") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"27F6C26BB7304972BC5C5B825ACC3771") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"46AB5D56";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"27F6C26BB7304972BC5C5B825ACC3771") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 673 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"46AB5D56") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BC330AD4557A66A7CE46C979D8527CD3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"46AB5D56";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BC330AD4557A66A7CE46C979D8527CD3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 674 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"46AB5D56") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D08B8AE0E2CCF649BE7669D5CC7A1536") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"46AB5D56";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D08B8AE0E2CCF649BE7669D5CC7A1536") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 675 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"46AB5D56") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8FEF2799FFE88D7E9B1A02956B1262F3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"46AB5D56";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8FEF2799FFE88D7E9B1A02956B1262F3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 676 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"46AB5D56") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C9AB549BE3CA27BB01BA35390530E605") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"46AB5D56";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C9AB549BE3CA27BB01BA35390530E605") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 677 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"46AB5D56") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6C8D68622A8AB46F0AEFFB5AE313D781") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"46AB5D56";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6C8D68622A8AB46F0AEFFB5AE313D781") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 678 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"46AB5D56") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"76FC8965F00103BAF092BA70682A28BD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"46AB5D56";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"76FC8965F00103BAF092BA70682A28BD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 679 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"46AB5D56") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"071D14D26938AF8988698F759B8D5F3C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"46AB5D56";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"071D14D26938AF8988698F759B8D5F3C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 680 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"46AB5D56") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CD5098CCC193D962F8DDAC319AA82E49") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"46AB5D56";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CD5098CCC193D962F8DDAC319AA82E49") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 681 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"46AB5D56") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"45D1629F38A9DBE1608E58FF415CF118") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"46AB5D56";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"45D1629F38A9DBE1608E58FF415CF118") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 682 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"46AB5D56") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"598F0287DE5430B6BFF44B9D4AC547EB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"46AB5D56";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"598F0287DE5430B6BFF44B9D4AC547EB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 683 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"46AB5D56") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A859303BD83EAB6F25486322C7D44610") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"46AB5D56";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A859303BD83EAB6F25486322C7D44610") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 684 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"46AB5D56") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A72717463342458E6650F296BB2AC535") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"46AB5D56";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A72717463342458E6650F296BB2AC535") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 685 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"46AB5D56") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"418CA63AAAE26667B6D436F77DB3473B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"46AB5D56";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"418CA63AAAE26667B6D436F77DB3473B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 686 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"46AB5D56") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"832E95F9362829FF3EC5A89C4A690C0B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"46AB5D56";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"832E95F9362829FF3EC5A89C4A690C0B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 687 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"46AB5D56") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"27E245D7CCCC8F0698D90CE89EAB3E88") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"46AB5D56";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"27E245D7CCCC8F0698D90CE89EAB3E88") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 688 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"46AB5D56") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C58D77CA178D7C069256E09B1CB607DE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"46AB5D56";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C58D77CA178D7C069256E09B1CB607DE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 689 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"46AB5D56") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B9AB2EDC37469C3FBCC78547384A3CEA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"46AB5D56";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B9AB2EDC37469C3FBCC78547384A3CEA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 690 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"46AB5D56") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AE2C6B3ABCC85FE7589D21D10F86FD04") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"46AB5D56";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AE2C6B3ABCC85FE7589D21D10F86FD04") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 691 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"46AB5D56") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5602A0602841F7BF3BD3AC329A6D4D96") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"46AB5D56";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5602A0602841F7BF3BD3AC329A6D4D96") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 692 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"46AB5D56") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"02362D05068A3B0C6D929C299DC604FA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"46AB5D56";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"02362D05068A3B0C6D929C299DC604FA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 693 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"46AB5D56") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E45B97BB72E346AC9A5CAF2A3899E177") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"46AB5D56";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-3)) = x"10111213") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E45B97BB72E346AC9A5CAF2A3899E177") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 694 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"46AB5D5674") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7CD0AD142A546E1C399ED92972EA5A66") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"46AB5D5674";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7CD0AD142A546E1C399ED92972EA5A66") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 695 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"46AB5D5674") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8A5C2D414E4BB653DE9453F1A4AD8945") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"46AB5D5674";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8A5C2D414E4BB653DE9453F1A4AD8945") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 696 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"46AB5D5674") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0719A0D604FFF3D1A33E32E428BDAE47") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"46AB5D5674";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0719A0D604FFF3D1A33E32E428BDAE47") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 697 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"46AB5D5674") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D3F4943A5FEE596A0238C89F0CA61ED6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"46AB5D5674";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D3F4943A5FEE596A0238C89F0CA61ED6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 698 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"46AB5D5674") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"42B98C0096725867E59DF0DF9DD1D239") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"46AB5D5674";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"42B98C0096725867E59DF0DF9DD1D239") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 699 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"46AB5D5674") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"600BF7F2EB777FC2B39B1DD464F6B4D6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"46AB5D5674";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"600BF7F2EB777FC2B39B1DD464F6B4D6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 700 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"46AB5D5674") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F57A0A1C366BB163158874965B072695") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"46AB5D5674";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F57A0A1C366BB163158874965B072695") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 701 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"46AB5D5674") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"44EA0604F02480D84A7B8BBBB1A0A98D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"46AB5D5674";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"44EA0604F02480D84A7B8BBBB1A0A98D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 702 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"46AB5D5674") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F7E2C6E899609F398D9DE7B2A56F035F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"46AB5D5674";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F7E2C6E899609F398D9DE7B2A56F035F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 703 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"46AB5D5674") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2BEEAD60817FDE6EE96A70BE0788F3C6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"46AB5D5674";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2BEEAD60817FDE6EE96A70BE0788F3C6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 704 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"46AB5D5674") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9BF6763A57D8D72FA850B7BC986469FD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"46AB5D5674";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9BF6763A57D8D72FA850B7BC986469FD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 705 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"46AB5D5674") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E4F99F6EAB9A280C23C5DB34F9174299") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"46AB5D5674";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E4F99F6EAB9A280C23C5DB34F9174299") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 706 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"46AB5D5674") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7F3C57D149D007D951DF49CF7B89093B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"46AB5D5674";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7F3C57D149D007D951DF49CF7B89093B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 707 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"46AB5D5674") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1384D7E5FE66973721EFE9636FA160DE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"46AB5D5674";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1384D7E5FE66973721EFE9636FA160DE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 708 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"46AB5D5674") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4CE07A9CE342EC0004838223C8C9171B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"46AB5D5674";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4CE07A9CE342EC0004838223C8C9171B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 709 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"46AB5D5674") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0AA4099EFF6046C59E23B58FA6EB93ED") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"46AB5D5674";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0AA4099EFF6046C59E23B58FA6EB93ED") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 710 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"46AB5D5674") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AF8235673620D51195767BEC40C8A269") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"46AB5D5674";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AF8235673620D51195767BEC40C8A269") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 711 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"46AB5D5674") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B5F3D460ECAB62C46F0B3AC6CBF15D55") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"46AB5D5674";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B5F3D460ECAB62C46F0B3AC6CBF15D55") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 712 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"46AB5D5674") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C41249D77592CEF717F00FC338562AD4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"46AB5D5674";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C41249D77592CEF717F00FC338562AD4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 713 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"46AB5D5674") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0E5FC5C9DD39B81C67442C8739735BA1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"46AB5D5674";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0E5FC5C9DD39B81C67442C8739735BA1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 714 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"46AB5D5674") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"86DE3F9A2403BA9FFF17D849E28784F0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"46AB5D5674";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"86DE3F9A2403BA9FFF17D849E28784F0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 715 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"46AB5D5674") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9A805F82C2FE51C8206DCB2BE91E3203") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"46AB5D5674";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9A805F82C2FE51C8206DCB2BE91E3203") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 716 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"46AB5D5674") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6B566D3EC494CA11BAD1E394640F33F8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"46AB5D5674";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6B566D3EC494CA11BAD1E394640F33F8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 717 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"46AB5D5674") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"64284A432FE824F0F9C9722018F1B0DD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"46AB5D5674";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"64284A432FE824F0F9C9722018F1B0DD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 718 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"46AB5D5674") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8283FB3FB6480719294DB641DE6832D3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"46AB5D5674";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8283FB3FB6480719294DB641DE6832D3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 719 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"46AB5D5674") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4021C8FC2A824881A15C282AE9B279E3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"46AB5D5674";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4021C8FC2A824881A15C282AE9B279E3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 720 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"46AB5D5674") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E4ED18D2D066EE7807408C5E3D704B60") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"46AB5D5674";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E4ED18D2D066EE7807408C5E3D704B60") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 721 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"46AB5D5674") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"06822ACF0B271D780DCF602DBF6D7236") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"46AB5D5674";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"06822ACF0B271D780DCF602DBF6D7236") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 722 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"46AB5D5674") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7AA473D92BECFD41235E05F19B914902") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"46AB5D5674";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7AA473D92BECFD41235E05F19B914902") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 723 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"46AB5D5674") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6D23363FA0623E99C704A167AC5D88EC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"46AB5D5674";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6D23363FA0623E99C704A167AC5D88EC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 724 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"46AB5D5674") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"950DFD6534EB96C1A44A2C8439B6387E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"46AB5D5674";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"950DFD6534EB96C1A44A2C8439B6387E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 725 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"46AB5D5674") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C13970001A205A72F20B1C9F3E1D7112") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"46AB5D5674";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C13970001A205A72F20B1C9F3E1D7112") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 726 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"46AB5D5674") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2754CABE6E4927D205C52F9C9B42949F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"46AB5D5674";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-4)) = x"1011121314") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2754CABE6E4927D205C52F9C9B42949F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 727 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"46AB5D56747C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8CEF300691D56A1B047F25594D791661") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"46AB5D56747C";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8CEF300691D56A1B047F25594D791661") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 728 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"46AB5D56747C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7A63B053F5CAB254E375AF819B3EC542") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"46AB5D56747C";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7A63B053F5CAB254E375AF819B3EC542") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 729 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"46AB5D56747C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F7263DC4BF7EF7D69EDFCE94172EE240") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"46AB5D56747C";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F7263DC4BF7EF7D69EDFCE94172EE240") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 730 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"46AB5D56747C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"23CB0928E46F5D6D3FD934EF333552D1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"46AB5D56747C";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"23CB0928E46F5D6D3FD934EF333552D1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 731 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"46AB5D56747C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B28611122DF35C60D87C0CAFA2429E3E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"46AB5D56747C";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B28611122DF35C60D87C0CAFA2429E3E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 732 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"46AB5D56747C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"90346AE050F67BC58E7AE1A45B65F8D1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"46AB5D56747C";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"90346AE050F67BC58E7AE1A45B65F8D1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 733 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"46AB5D56747C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0545970E8DEAB564286988E664946A92") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"46AB5D56747C";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0545970E8DEAB564286988E664946A92") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 734 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"46AB5D56747C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B4D59B164BA584DF779A77CB8E33E58A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"46AB5D56747C";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B4D59B164BA584DF779A77CB8E33E58A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 735 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"46AB5D56747C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"07DD5BFA22E19B3EB07C1BC29AFC4F58") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"46AB5D56747C";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"07DD5BFA22E19B3EB07C1BC29AFC4F58") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 736 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"46AB5D56747C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DBD130723AFEDA69D48B8CCE381BBFC1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"46AB5D56747C";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DBD130723AFEDA69D48B8CCE381BBFC1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 737 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"46AB5D56747C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6BC9EB28EC59D32895B14BCCA7F725FA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"46AB5D56747C";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6BC9EB28EC59D32895B14BCCA7F725FA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 738 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"46AB5D56747C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"14C6027C101B2C0B1E242744C6840E9E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"46AB5D56747C";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"14C6027C101B2C0B1E242744C6840E9E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 739 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"46AB5D56747C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8F03CAC3F25103DE6C3EB5BF441A453C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"46AB5D56747C";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8F03CAC3F25103DE6C3EB5BF441A453C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 740 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"46AB5D56747C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E3BB4AF745E793301C0E151350322CD9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"46AB5D56747C";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E3BB4AF745E793301C0E151350322CD9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 741 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"46AB5D56747C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BCDFE78E58C3E80739627E53F75A5B1C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"46AB5D56747C";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BCDFE78E58C3E80739627E53F75A5B1C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 742 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"46AB5D56747C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FA9B948C44E142C2A3C249FF9978DFEA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"46AB5D56747C";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FA9B948C44E142C2A3C249FF9978DFEA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 743 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"46AB5D56747C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5FBDA8758DA1D116A897879C7F5BEE6E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"46AB5D56747C";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5FBDA8758DA1D116A897879C7F5BEE6E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 744 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"46AB5D56747C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"45CC4972572A66C352EAC6B6F4621152") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"46AB5D56747C";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"45CC4972572A66C352EAC6B6F4621152") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 745 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"46AB5D56747C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"342DD4C5CE13CAF02A11F3B307C566D3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"46AB5D56747C";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"342DD4C5CE13CAF02A11F3B307C566D3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 746 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"46AB5D56747C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FE6058DB66B8BC1B5AA5D0F706E017A6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"46AB5D56747C";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FE6058DB66B8BC1B5AA5D0F706E017A6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 747 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"46AB5D56747C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"76E1A2889F82BE98C2F62439DD14C8F7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"46AB5D56747C";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"76E1A2889F82BE98C2F62439DD14C8F7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 748 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"46AB5D56747C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6ABFC290797F55CF1D8C375BD68D7E04") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"46AB5D56747C";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6ABFC290797F55CF1D8C375BD68D7E04") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 749 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"46AB5D56747C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9B69F02C7F15CE1687301FE45B9C7FFF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"46AB5D56747C";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9B69F02C7F15CE1687301FE45B9C7FFF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 750 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"46AB5D56747C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9417D751946920F7C4288E502762FCDA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"46AB5D56747C";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9417D751946920F7C4288E502762FCDA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 751 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"46AB5D56747C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"72BC662D0DC9031E14AC4A31E1FB7ED4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"46AB5D56747C";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"72BC662D0DC9031E14AC4A31E1FB7ED4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 752 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"46AB5D56747C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B01E55EE91034C869CBDD45AD62135E4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"46AB5D56747C";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B01E55EE91034C869CBDD45AD62135E4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 753 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"46AB5D56747C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"14D285C06BE7EA7F3AA1702E02E30767") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"46AB5D56747C";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"14D285C06BE7EA7F3AA1702E02E30767") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 754 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"46AB5D56747C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F6BDB7DDB0A6197F302E9C5D80FE3E31") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"46AB5D56747C";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F6BDB7DDB0A6197F302E9C5D80FE3E31") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 755 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"46AB5D56747C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8A9BEECB906DF9461EBFF981A4020505") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"46AB5D56747C";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8A9BEECB906DF9461EBFF981A4020505") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 756 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"46AB5D56747C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9D1CAB2D1BE33A9EFAE55D1793CEC4EB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"46AB5D56747C";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9D1CAB2D1BE33A9EFAE55D1793CEC4EB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 757 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"46AB5D56747C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"653260778F6A92C699ABD0F406257479") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"46AB5D56747C";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"653260778F6A92C699ABD0F406257479") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 758 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"46AB5D56747C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3106ED12A1A15E75CFEAE0EF018E3D15") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"46AB5D56747C";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3106ED12A1A15E75CFEAE0EF018E3D15") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 759 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"46AB5D56747C") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D76B57ACD5C823D53824D3ECA4D1D898") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"46AB5D56747C";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-5)) = x"101112131415") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D76B57ACD5C823D53824D3ECA4D1D898") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 760 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"46AB5D56747C33") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0BAE8A9FA9565D0AB9158E038160C107") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"46AB5D56747C33";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0BAE8A9FA9565D0AB9158E038160C107") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 761 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"46AB5D56747C33") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FD220ACACD4985455E1F04DB57271224") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"46AB5D56747C33";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FD220ACACD4985455E1F04DB57271224") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 762 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"46AB5D56747C33") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7067875D87FDC0C723B565CEDB373526") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"46AB5D56747C33";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7067875D87FDC0C723B565CEDB373526") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 763 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"46AB5D56747C33") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A48AB3B1DCEC6A7C82B39FB5FF2C85B7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"46AB5D56747C33";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A48AB3B1DCEC6A7C82B39FB5FF2C85B7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 764 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"46AB5D56747C33") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"35C7AB8B15706B716516A7F56E5B4958") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"46AB5D56747C33";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"35C7AB8B15706B716516A7F56E5B4958") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 765 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"46AB5D56747C33") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1775D07968754CD433104AFE977C2FB7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"46AB5D56747C33";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1775D07968754CD433104AFE977C2FB7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 766 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"46AB5D56747C33") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"82042D97B5698275950323BCA88DBDF4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"46AB5D56747C33";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"82042D97B5698275950323BCA88DBDF4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 767 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"46AB5D56747C33") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3394218F7326B3CECAF0DC91422A32EC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"46AB5D56747C33";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3394218F7326B3CECAF0DC91422A32EC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 768 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"46AB5D56747C33") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"809CE1631A62AC2F0D16B09856E5983E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"46AB5D56747C33";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"809CE1631A62AC2F0D16B09856E5983E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 769 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"46AB5D56747C33") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5C908AEB027DED7869E12794F40268A7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"46AB5D56747C33";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5C908AEB027DED7869E12794F40268A7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 770 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"46AB5D56747C33") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EC8851B1D4DAE43928DBE0966BEEF29C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"46AB5D56747C33";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EC8851B1D4DAE43928DBE0966BEEF29C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 771 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"46AB5D56747C33") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9387B8E528981B1AA34E8C1E0A9DD9F8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"46AB5D56747C33";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9387B8E528981B1AA34E8C1E0A9DD9F8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 772 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"46AB5D56747C33") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0842705ACAD234CFD1541EE58803925A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"46AB5D56747C33";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0842705ACAD234CFD1541EE58803925A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 773 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"46AB5D56747C33") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"64FAF06E7D64A421A164BE499C2BFBBF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"46AB5D56747C33";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"64FAF06E7D64A421A164BE499C2BFBBF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 774 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"46AB5D56747C33") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3B9E5D176040DF168408D5093B438C7A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"46AB5D56747C33";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3B9E5D176040DF168408D5093B438C7A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 775 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"46AB5D56747C33") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7DDA2E157C6275D31EA8E2A55561088C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"46AB5D56747C33";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7DDA2E157C6275D31EA8E2A55561088C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 776 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"46AB5D56747C33") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D8FC12ECB522E60715FD2CC6B3423908") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"46AB5D56747C33";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D8FC12ECB522E60715FD2CC6B3423908") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 777 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"46AB5D56747C33") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C28DF3EB6FA951D2EF806DEC387BC634") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"46AB5D56747C33";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C28DF3EB6FA951D2EF806DEC387BC634") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 778 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"46AB5D56747C33") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B36C6E5CF690FDE1977B58E9CBDCB1B5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"46AB5D56747C33";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B36C6E5CF690FDE1977B58E9CBDCB1B5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 779 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"46AB5D56747C33") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7921E2425E3B8B0AE7CF7BADCAF9C0C0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"46AB5D56747C33";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7921E2425E3B8B0AE7CF7BADCAF9C0C0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 780 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"46AB5D56747C33") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F1A01811A70189897F9C8F63110D1F91") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"46AB5D56747C33";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F1A01811A70189897F9C8F63110D1F91") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 781 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"46AB5D56747C33") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EDFE780941FC62DEA0E69C011A94A962") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"46AB5D56747C33";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EDFE780941FC62DEA0E69C011A94A962") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 782 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"46AB5D56747C33") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1C284AB54796F9073A5AB4BE9785A899") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"46AB5D56747C33";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1C284AB54796F9073A5AB4BE9785A899") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 783 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"46AB5D56747C33") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"13566DC8ACEA17E67942250AEB7B2BBC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"46AB5D56747C33";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"13566DC8ACEA17E67942250AEB7B2BBC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 784 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"46AB5D56747C33") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F5FDDCB4354A340FA9C6E16B2DE2A9B2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"46AB5D56747C33";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F5FDDCB4354A340FA9C6E16B2DE2A9B2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 785 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"46AB5D56747C33") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"375FEF77A9807B9721D77F001A38E282") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"46AB5D56747C33";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"375FEF77A9807B9721D77F001A38E282") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 786 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"46AB5D56747C33") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"93933F595364DD6E87CBDB74CEFAD001") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"46AB5D56747C33";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"93933F595364DD6E87CBDB74CEFAD001") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 787 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"46AB5D56747C33") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"71FC0D4488252E6E8D4437074CE7E957") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"46AB5D56747C33";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"71FC0D4488252E6E8D4437074CE7E957") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 788 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"46AB5D56747C33") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0DDA5452A8EECE57A3D552DB681BD263") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"46AB5D56747C33";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0DDA5452A8EECE57A3D552DB681BD263") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 789 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"46AB5D56747C33") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1A5D11B423600D8F478FF64D5FD7138D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"46AB5D56747C33";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1A5D11B423600D8F478FF64D5FD7138D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 790 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"46AB5D56747C33") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E273DAEEB7E9A5D724C17BAECA3CA31F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"46AB5D56747C33";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E273DAEEB7E9A5D724C17BAECA3CA31F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 791 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"46AB5D56747C33") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B647578B9922696472804BB5CD97EA73") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"46AB5D56747C33";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B647578B9922696472804BB5CD97EA73") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 792 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"46AB5D56747C33") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"502AED35ED4B14C4854E78B668C80FFE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"46AB5D56747C33";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-6)) = x"10111213141516") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"502AED35ED4B14C4854E78B668C80FFE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 793 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"46AB5D56747C33F9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"386E25E16BF47889C037CE63DD4FCF33") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"46AB5D56747C33F9";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"386E25E16BF47889C037CE63DD4FCF33") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 794 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"46AB5D56747C33F9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CEE2A5B40FEBA0C6273D44BB0B081C10") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"46AB5D56747C33F9";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CEE2A5B40FEBA0C6273D44BB0B081C10") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 795 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"46AB5D56747C33F9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"43A72823455FE5445A9725AE87183B12") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"46AB5D56747C33F9";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"43A72823455FE5445A9725AE87183B12") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 796 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"46AB5D56747C33F9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"974A1CCF1E4E4FFFFB91DFD5A3038B83") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"46AB5D56747C33F9";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"974A1CCF1E4E4FFFFB91DFD5A3038B83") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 797 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"46AB5D56747C33F9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"060704F5D7D24EF21C34E7953274476C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"46AB5D56747C33F9";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"060704F5D7D24EF21C34E7953274476C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 798 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"46AB5D56747C33F9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"24B57F07AAD769574A320A9ECB532183") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"46AB5D56747C33F9";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"24B57F07AAD769574A320A9ECB532183") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 799 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"46AB5D56747C33F9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B1C482E977CBA7F6EC2163DCF4A2B3C0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"46AB5D56747C33F9";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B1C482E977CBA7F6EC2163DCF4A2B3C0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 800 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"46AB5D56747C33F9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"00548EF1B184964DB3D29CF11E053CD8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"46AB5D56747C33F9";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"00548EF1B184964DB3D29CF11E053CD8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 801 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"46AB5D56747C33F9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B35C4E1DD8C089AC7434F0F80ACA960A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"46AB5D56747C33F9";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B35C4E1DD8C089AC7434F0F80ACA960A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 802 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"46AB5D56747C33F9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6F502595C0DFC8FB10C367F4A82D6693") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"46AB5D56747C33F9";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6F502595C0DFC8FB10C367F4A82D6693") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 803 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"46AB5D56747C33F9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DF48FECF1678C1BA51F9A0F637C1FCA8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"46AB5D56747C33F9";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DF48FECF1678C1BA51F9A0F637C1FCA8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 804 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"46AB5D56747C33F9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A047179BEA3A3E99DA6CCC7E56B2D7CC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"46AB5D56747C33F9";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A047179BEA3A3E99DA6CCC7E56B2D7CC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 805 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"46AB5D56747C33F9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3B82DF240870114CA8765E85D42C9C6E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"46AB5D56747C33F9";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3B82DF240870114CA8765E85D42C9C6E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 806 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"46AB5D56747C33F9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"573A5F10BFC681A2D846FE29C004F58B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"46AB5D56747C33F9";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"573A5F10BFC681A2D846FE29C004F58B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 807 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"46AB5D56747C33F9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"085EF269A2E2FA95FD2A9569676C824E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"46AB5D56747C33F9";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"085EF269A2E2FA95FD2A9569676C824E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 808 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"46AB5D56747C33F9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4E1A816BBEC05050678AA2C5094E06B8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"46AB5D56747C33F9";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4E1A816BBEC05050678AA2C5094E06B8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 809 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"46AB5D56747C33F9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EB3CBD927780C3846CDF6CA6EF6D373C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"46AB5D56747C33F9";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EB3CBD927780C3846CDF6CA6EF6D373C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 810 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"46AB5D56747C33F9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F14D5C95AD0B745196A22D8C6454C800") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"46AB5D56747C33F9";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F14D5C95AD0B745196A22D8C6454C800") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 811 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"46AB5D56747C33F9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"80ACC1223432D862EE59188997F3BF81") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"46AB5D56747C33F9";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"80ACC1223432D862EE59188997F3BF81") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 812 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"46AB5D56747C33F9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4AE14D3C9C99AE899EED3BCD96D6CEF4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"46AB5D56747C33F9";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4AE14D3C9C99AE899EED3BCD96D6CEF4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 813 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"46AB5D56747C33F9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C260B76F65A3AC0A06BECF034D2211A5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"46AB5D56747C33F9";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C260B76F65A3AC0A06BECF034D2211A5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 814 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"46AB5D56747C33F9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DE3ED777835E475DD9C4DC6146BBA756") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"46AB5D56747C33F9";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DE3ED777835E475DD9C4DC6146BBA756") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 815 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"46AB5D56747C33F9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2FE8E5CB8534DC844378F4DECBAAA6AD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"46AB5D56747C33F9";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2FE8E5CB8534DC844378F4DECBAAA6AD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 816 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"46AB5D56747C33F9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2096C2B66E4832650060656AB7542588") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"46AB5D56747C33F9";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2096C2B66E4832650060656AB7542588") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 817 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"46AB5D56747C33F9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C63D73CAF7E8118CD0E4A10B71CDA786") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"46AB5D56747C33F9";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C63D73CAF7E8118CD0E4A10B71CDA786") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 818 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"46AB5D56747C33F9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"049F40096B225E1458F53F604617ECB6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"46AB5D56747C33F9";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"049F40096B225E1458F53F604617ECB6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 819 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"46AB5D56747C33F9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A053902791C6F8EDFEE99B1492D5DE35") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"46AB5D56747C33F9";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A053902791C6F8EDFEE99B1492D5DE35") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 820 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"46AB5D56747C33F9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"423CA23A4A870BEDF466776710C8E763") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"46AB5D56747C33F9";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"423CA23A4A870BEDF466776710C8E763") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 821 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"46AB5D56747C33F9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3E1AFB2C6A4CEBD4DAF712BB3434DC57") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"46AB5D56747C33F9";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3E1AFB2C6A4CEBD4DAF712BB3434DC57") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 822 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"46AB5D56747C33F9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"299DBECAE1C2280C3EADB62D03F81DB9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"46AB5D56747C33F9";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"299DBECAE1C2280C3EADB62D03F81DB9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 823 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"46AB5D56747C33F9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D1B37590754B80545DE33BCE9613AD2B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"46AB5D56747C33F9";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D1B37590754B80545DE33BCE9613AD2B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 824 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"46AB5D56747C33F9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8587F8F55B804CE70BA20BD591B8E447") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"46AB5D56747C33F9";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8587F8F55B804CE70BA20BD591B8E447") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 825 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"46AB5D56747C33F9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"63EA424B2FE93147FC6C38D634E701CA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"46AB5D56747C33F9";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-7)) = x"1011121314151617") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"63EA424B2FE93147FC6C38D634E701CA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 826 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"46AB5D56747C33F905") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0122F7023366642DC6A67804E3304605") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"46AB5D56747C33F905";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0122F7023366642DC6A67804E3304605") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 827 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"46AB5D56747C33F905") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F7AE77575779BC6221ACF2DC35779526") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"46AB5D56747C33F905";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F7AE77575779BC6221ACF2DC35779526") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 828 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"46AB5D56747C33F905") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7AEBFAC01DCDF9E05C0693C9B967B224") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"46AB5D56747C33F905";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7AEBFAC01DCDF9E05C0693C9B967B224") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 829 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"46AB5D56747C33F905") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AE06CE2C46DC535BFD0069B29D7C02B5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"46AB5D56747C33F905";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AE06CE2C46DC535BFD0069B29D7C02B5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 830 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"46AB5D56747C33F905") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3F4BD6168F4052561AA551F20C0BCE5A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"46AB5D56747C33F905";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3F4BD6168F4052561AA551F20C0BCE5A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 831 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"46AB5D56747C33F905") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1DF9ADE4F24575F34CA3BCF9F52CA8B5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"46AB5D56747C33F905";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1DF9ADE4F24575F34CA3BCF9F52CA8B5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 832 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"46AB5D56747C33F905") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8888500A2F59BB52EAB0D5BBCADD3AF6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"46AB5D56747C33F905";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8888500A2F59BB52EAB0D5BBCADD3AF6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 833 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"46AB5D56747C33F905") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"39185C12E9168AE9B5432A96207AB5EE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"46AB5D56747C33F905";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"39185C12E9168AE9B5432A96207AB5EE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 834 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"46AB5D56747C33F905") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8A109CFE8052950872A5469F34B51F3C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"46AB5D56747C33F905";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8A109CFE8052950872A5469F34B51F3C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 835 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"46AB5D56747C33F905") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"561CF776984DD45F1652D1939652EFA5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"46AB5D56747C33F905";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"561CF776984DD45F1652D1939652EFA5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 836 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"46AB5D56747C33F905") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E6042C2C4EEADD1E5768169109BE759E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"46AB5D56747C33F905";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E6042C2C4EEADD1E5768169109BE759E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 837 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"46AB5D56747C33F905") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"990BC578B2A8223DDCFD7A1968CD5EFA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"46AB5D56747C33F905";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"990BC578B2A8223DDCFD7A1968CD5EFA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 838 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"46AB5D56747C33F905") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"02CE0DC750E20DE8AEE7E8E2EA531558") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"46AB5D56747C33F905";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"02CE0DC750E20DE8AEE7E8E2EA531558") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 839 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"46AB5D56747C33F905") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6E768DF3E7549D06DED7484EFE7B7CBD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"46AB5D56747C33F905";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6E768DF3E7549D06DED7484EFE7B7CBD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 840 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"46AB5D56747C33F905") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3112208AFA70E631FBBB230E59130B78") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"46AB5D56747C33F905";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3112208AFA70E631FBBB230E59130B78") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 841 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"46AB5D56747C33F905") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"77565388E6524CF4611B14A237318F8E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"46AB5D56747C33F905";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"77565388E6524CF4611B14A237318F8E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 842 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"46AB5D56747C33F905") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D2706F712F12DF206A4EDAC1D112BE0A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"46AB5D56747C33F905";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D2706F712F12DF206A4EDAC1D112BE0A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 843 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"46AB5D56747C33F905") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C8018E76F59968F590339BEB5A2B4136") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"46AB5D56747C33F905";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C8018E76F59968F590339BEB5A2B4136") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 844 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"46AB5D56747C33F905") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B9E013C16CA0C4C6E8C8AEEEA98C36B7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"46AB5D56747C33F905";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B9E013C16CA0C4C6E8C8AEEEA98C36B7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 845 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"46AB5D56747C33F905") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"73AD9FDFC40BB22D987C8DAAA8A947C2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"46AB5D56747C33F905";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"73AD9FDFC40BB22D987C8DAAA8A947C2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 846 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"46AB5D56747C33F905") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FB2C658C3D31B0AE002F7964735D9893") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"46AB5D56747C33F905";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FB2C658C3D31B0AE002F7964735D9893") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 847 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"46AB5D56747C33F905") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E7720594DBCC5BF9DF556A0678C42E60") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"46AB5D56747C33F905";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E7720594DBCC5BF9DF556A0678C42E60") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 848 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"46AB5D56747C33F905") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"16A43728DDA6C02045E942B9F5D52F9B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"46AB5D56747C33F905";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"16A43728DDA6C02045E942B9F5D52F9B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 849 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"46AB5D56747C33F905") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"19DA105536DA2EC106F1D30D892BACBE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"46AB5D56747C33F905";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"19DA105536DA2EC106F1D30D892BACBE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 850 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"46AB5D56747C33F905") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FF71A129AF7A0D28D675176C4FB22EB0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"46AB5D56747C33F905";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FF71A129AF7A0D28D675176C4FB22EB0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 851 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"46AB5D56747C33F905") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3DD392EA33B042B05E64890778686580") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"46AB5D56747C33F905";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3DD392EA33B042B05E64890778686580") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 852 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"46AB5D56747C33F905") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"991F42C4C954E449F8782D73ACAA5703") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"46AB5D56747C33F905";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"991F42C4C954E449F8782D73ACAA5703") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 853 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"46AB5D56747C33F905") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7B7070D912151749F2F7C1002EB76E55") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"46AB5D56747C33F905";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7B7070D912151749F2F7C1002EB76E55") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 854 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"46AB5D56747C33F905") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"075629CF32DEF770DC66A4DC0A4B5561") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"46AB5D56747C33F905";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"075629CF32DEF770DC66A4DC0A4B5561") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 855 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"46AB5D56747C33F905") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"10D16C29B95034A8383C004A3D87948F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"46AB5D56747C33F905";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"10D16C29B95034A8383C004A3D87948F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 856 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"46AB5D56747C33F905") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E8FFA7732DD99CF05B728DA9A86C241D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"46AB5D56747C33F905";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E8FFA7732DD99CF05B728DA9A86C241D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 857 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"46AB5D56747C33F905") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BCCB2A16031250430D33BDB2AFC76D71") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"46AB5D56747C33F905";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BCCB2A16031250430D33BDB2AFC76D71") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 858 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"46AB5D56747C33F905") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5AA690A8777B2DE3FAFD8EB10A9888FC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"46AB5D56747C33F905";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-8)) = x"101112131415161718") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5AA690A8777B2DE3FAFD8EB10A9888FC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 859 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"46AB5D56747C33F90529") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EC667DBD737AA315D9E9B026038B6747") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"46AB5D56747C33F90529";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EC667DBD737AA315D9E9B026038B6747") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 860 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"46AB5D56747C33F90529") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1AEAFDE817657B5A3EE33AFED5CCB464") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"46AB5D56747C33F90529";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1AEAFDE817657B5A3EE33AFED5CCB464") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 861 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"46AB5D56747C33F90529") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"97AF707F5DD13ED843495BEB59DC9366") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"46AB5D56747C33F90529";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"97AF707F5DD13ED843495BEB59DC9366") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 862 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"46AB5D56747C33F90529") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4342449306C09463E24FA1907DC723F7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"46AB5D56747C33F90529";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4342449306C09463E24FA1907DC723F7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 863 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"46AB5D56747C33F90529") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D20F5CA9CF5C956E05EA99D0ECB0EF18") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"46AB5D56747C33F90529";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D20F5CA9CF5C956E05EA99D0ECB0EF18") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 864 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"46AB5D56747C33F90529") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F0BD275BB259B2CB53EC74DB159789F7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"46AB5D56747C33F90529";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F0BD275BB259B2CB53EC74DB159789F7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 865 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"46AB5D56747C33F90529") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"65CCDAB56F457C6AF5FF1D992A661BB4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"46AB5D56747C33F90529";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"65CCDAB56F457C6AF5FF1D992A661BB4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 866 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"46AB5D56747C33F90529") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D45CD6ADA90A4DD1AA0CE2B4C0C194AC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"46AB5D56747C33F90529";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D45CD6ADA90A4DD1AA0CE2B4C0C194AC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 867 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"46AB5D56747C33F90529") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"67541641C04E52306DEA8EBDD40E3E7E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"46AB5D56747C33F90529";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"67541641C04E52306DEA8EBDD40E3E7E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 868 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"46AB5D56747C33F90529") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BB587DC9D8511367091D19B176E9CEE7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"46AB5D56747C33F90529";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BB587DC9D8511367091D19B176E9CEE7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 869 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"46AB5D56747C33F90529") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0B40A6930EF61A264827DEB3E90554DC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"46AB5D56747C33F90529";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0B40A6930EF61A264827DEB3E90554DC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 870 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"46AB5D56747C33F90529") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"744F4FC7F2B4E505C3B2B23B88767FB8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"46AB5D56747C33F90529";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"744F4FC7F2B4E505C3B2B23B88767FB8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 871 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"46AB5D56747C33F90529") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EF8A877810FECAD0B1A820C00AE8341A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"46AB5D56747C33F90529";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EF8A877810FECAD0B1A820C00AE8341A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 872 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"46AB5D56747C33F90529") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8332074CA7485A3EC198806C1EC05DFF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"46AB5D56747C33F90529";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8332074CA7485A3EC198806C1EC05DFF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 873 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"46AB5D56747C33F90529") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DC56AA35BA6C2109E4F4EB2CB9A82A3A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"46AB5D56747C33F90529";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DC56AA35BA6C2109E4F4EB2CB9A82A3A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 874 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"46AB5D56747C33F90529") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9A12D937A64E8BCC7E54DC80D78AAECC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"46AB5D56747C33F90529";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9A12D937A64E8BCC7E54DC80D78AAECC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 875 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"46AB5D56747C33F90529") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3F34E5CE6F0E1818750112E331A99F48") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"46AB5D56747C33F90529";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3F34E5CE6F0E1818750112E331A99F48") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 876 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"46AB5D56747C33F90529") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"254504C9B585AFCD8F7C53C9BA906074") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"46AB5D56747C33F90529";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"254504C9B585AFCD8F7C53C9BA906074") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 877 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"46AB5D56747C33F90529") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"54A4997E2CBC03FEF78766CC493717F5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"46AB5D56747C33F90529";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"54A4997E2CBC03FEF78766CC493717F5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 878 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"46AB5D56747C33F90529") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9EE91560841775158733458848126680") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"46AB5D56747C33F90529";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9EE91560841775158733458848126680") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 879 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"46AB5D56747C33F90529") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1668EF337D2D77961F60B14693E6B9D1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"46AB5D56747C33F90529";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1668EF337D2D77961F60B14693E6B9D1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 880 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"46AB5D56747C33F90529") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0A368F2B9BD09CC1C01AA224987F0F22") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"46AB5D56747C33F90529";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0A368F2B9BD09CC1C01AA224987F0F22") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 881 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"46AB5D56747C33F90529") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FBE0BD979DBA07185AA68A9B156E0ED9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"46AB5D56747C33F90529";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FBE0BD979DBA07185AA68A9B156E0ED9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 882 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"46AB5D56747C33F90529") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F49E9AEA76C6E9F919BE1B2F69908DFC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"46AB5D56747C33F90529";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F49E9AEA76C6E9F919BE1B2F69908DFC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 883 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"46AB5D56747C33F90529") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"12352B96EF66CA10C93ADF4EAF090FF2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"46AB5D56747C33F90529";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"12352B96EF66CA10C93ADF4EAF090FF2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 884 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"46AB5D56747C33F90529") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D097185573AC8588412B412598D344C2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"46AB5D56747C33F90529";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D097185573AC8588412B412598D344C2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 885 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"46AB5D56747C33F90529") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"745BC87B89482371E737E5514C117641") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"46AB5D56747C33F90529";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"745BC87B89482371E737E5514C117641") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 886 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"46AB5D56747C33F90529") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9634FA665209D071EDB80922CE0C4F17") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"46AB5D56747C33F90529";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9634FA665209D071EDB80922CE0C4F17") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 887 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"46AB5D56747C33F90529") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EA12A37072C23048C3296CFEEAF07423") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"46AB5D56747C33F90529";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EA12A37072C23048C3296CFEEAF07423") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 888 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"46AB5D56747C33F90529") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FD95E696F94CF3902773C868DD3CB5CD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"46AB5D56747C33F90529";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FD95E696F94CF3902773C868DD3CB5CD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 889 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"46AB5D56747C33F90529") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"05BB2DCC6DC55BC8443D458B48D7055F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"46AB5D56747C33F90529";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"05BB2DCC6DC55BC8443D458B48D7055F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 890 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"46AB5D56747C33F90529") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"518FA0A9430E977B127C75904F7C4C33") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"46AB5D56747C33F90529";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"518FA0A9430E977B127C75904F7C4C33") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 891 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"46AB5D56747C33F90529") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B7E21A173767EADBE5B24693EA23A9BE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"46AB5D56747C33F90529";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-9)) = x"10111213141516171819") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B7E21A173767EADBE5B24693EA23A9BE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 892 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"46AB5D56747C33F9052911") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"16570F29C9FFB530F8512E916BD0B8D4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"46AB5D56747C33F9052911";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"16570F29C9FFB530F8512E916BD0B8D4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 893 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"46AB5D56747C33F9052911") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E0DB8F7CADE06D7F1F5BA449BD976BF7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"46AB5D56747C33F9052911";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E0DB8F7CADE06D7F1F5BA449BD976BF7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 894 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"46AB5D56747C33F9052911") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6D9E02EBE75428FD62F1C55C31874CF5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"46AB5D56747C33F9052911";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6D9E02EBE75428FD62F1C55C31874CF5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 895 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"46AB5D56747C33F9052911") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B9733607BC458246C3F73F27159CFC64") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"46AB5D56747C33F9052911";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B9733607BC458246C3F73F27159CFC64") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 896 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"46AB5D56747C33F9052911") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"283E2E3D75D9834B2452076784EB308B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"46AB5D56747C33F9052911";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"283E2E3D75D9834B2452076784EB308B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 897 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"46AB5D56747C33F9052911") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0A8C55CF08DCA4EE7254EA6C7DCC5664") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"46AB5D56747C33F9052911";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0A8C55CF08DCA4EE7254EA6C7DCC5664") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 898 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"46AB5D56747C33F9052911") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9FFDA821D5C06A4FD447832E423DC427") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"46AB5D56747C33F9052911";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9FFDA821D5C06A4FD447832E423DC427") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 899 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"46AB5D56747C33F9052911") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2E6DA439138F5BF48BB47C03A89A4B3F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"46AB5D56747C33F9052911";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2E6DA439138F5BF48BB47C03A89A4B3F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 900 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"46AB5D56747C33F9052911") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9D6564D57ACB44154C52100ABC55E1ED") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"46AB5D56747C33F9052911";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9D6564D57ACB44154C52100ABC55E1ED") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 901 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"46AB5D56747C33F9052911") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"41690F5D62D4054228A587061EB21174") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"46AB5D56747C33F9052911";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"41690F5D62D4054228A587061EB21174") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 902 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"46AB5D56747C33F9052911") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F171D407B4730C03699F4004815E8B4F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"46AB5D56747C33F9052911";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F171D407B4730C03699F4004815E8B4F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 903 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"46AB5D56747C33F9052911") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8E7E3D534831F320E20A2C8CE02DA02B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"46AB5D56747C33F9052911";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8E7E3D534831F320E20A2C8CE02DA02B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 904 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"46AB5D56747C33F9052911") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"15BBF5ECAA7BDCF59010BE7762B3EB89") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"46AB5D56747C33F9052911";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"15BBF5ECAA7BDCF59010BE7762B3EB89") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 905 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"46AB5D56747C33F9052911") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"790375D81DCD4C1BE0201EDB769B826C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"46AB5D56747C33F9052911";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"790375D81DCD4C1BE0201EDB769B826C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 906 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"46AB5D56747C33F9052911") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2667D8A100E9372CC54C759BD1F3F5A9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"46AB5D56747C33F9052911";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2667D8A100E9372CC54C759BD1F3F5A9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 907 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"46AB5D56747C33F9052911") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6023ABA31CCB9DE95FEC4237BFD1715F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"46AB5D56747C33F9052911";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6023ABA31CCB9DE95FEC4237BFD1715F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 908 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"46AB5D56747C33F9052911") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C505975AD58B0E3D54B98C5459F240DB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"46AB5D56747C33F9052911";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C505975AD58B0E3D54B98C5459F240DB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 909 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"46AB5D56747C33F9052911") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DF74765D0F00B9E8AEC4CD7ED2CBBFE7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"46AB5D56747C33F9052911";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DF74765D0F00B9E8AEC4CD7ED2CBBFE7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 910 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"46AB5D56747C33F9052911") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AE95EBEA963915DBD63FF87B216CC866") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"46AB5D56747C33F9052911";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AE95EBEA963915DBD63FF87B216CC866") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 911 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"46AB5D56747C33F9052911") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"64D867F43E926330A68BDB3F2049B913") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"46AB5D56747C33F9052911";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"64D867F43E926330A68BDB3F2049B913") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 912 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"46AB5D56747C33F9052911") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EC599DA7C7A861B33ED82FF1FBBD6642") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"46AB5D56747C33F9052911";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EC599DA7C7A861B33ED82FF1FBBD6642") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 913 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"46AB5D56747C33F9052911") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F007FDBF21558AE4E1A23C93F024D0B1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"46AB5D56747C33F9052911";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F007FDBF21558AE4E1A23C93F024D0B1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 914 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"46AB5D56747C33F9052911") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"01D1CF03273F113D7B1E142C7D35D14A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"46AB5D56747C33F9052911";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"01D1CF03273F113D7B1E142C7D35D14A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 915 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"46AB5D56747C33F9052911") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0EAFE87ECC43FFDC3806859801CB526F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"46AB5D56747C33F9052911";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0EAFE87ECC43FFDC3806859801CB526F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 916 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"46AB5D56747C33F9052911") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E804590255E3DC35E88241F9C752D061") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"46AB5D56747C33F9052911";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E804590255E3DC35E88241F9C752D061") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 917 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"46AB5D56747C33F9052911") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2AA66AC1C92993AD6093DF92F0889B51") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"46AB5D56747C33F9052911";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2AA66AC1C92993AD6093DF92F0889B51") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 918 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"46AB5D56747C33F9052911") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8E6ABAEF33CD3554C68F7BE6244AA9D2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"46AB5D56747C33F9052911";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8E6ABAEF33CD3554C68F7BE6244AA9D2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 919 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"46AB5D56747C33F9052911") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6C0588F2E88CC654CC009795A6579084") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"46AB5D56747C33F9052911";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6C0588F2E88CC654CC009795A6579084") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 920 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"46AB5D56747C33F9052911") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1023D1E4C847266DE291F24982ABABB0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"46AB5D56747C33F9052911";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1023D1E4C847266DE291F24982ABABB0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 921 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"46AB5D56747C33F9052911") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"07A4940243C9E5B506CB56DFB5676A5E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"46AB5D56747C33F9052911";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"07A4940243C9E5B506CB56DFB5676A5E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 922 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"46AB5D56747C33F9052911") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FF8A5F58D7404DED6585DB3C208CDACC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"46AB5D56747C33F9052911";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FF8A5F58D7404DED6585DB3C208CDACC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 923 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"46AB5D56747C33F9052911") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"ABBED23DF98B815E33C4EB27272793A0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"46AB5D56747C33F9052911";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"ABBED23DF98B815E33C4EB27272793A0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 924 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"46AB5D56747C33F9052911") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4DD368838DE2FCFEC40AD8248278762D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"46AB5D56747C33F9052911";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-10)) = x"101112131415161718191A") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4DD368838DE2FCFEC40AD8248278762D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 925 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"46AB5D56747C33F9052911BD") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"83537BC552DD0FB9D9EE96289F9FDC08") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"46AB5D56747C33F9052911BD";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"83537BC552DD0FB9D9EE96289F9FDC08") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 926 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"46AB5D56747C33F9052911BD") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"75DFFB9036C2D7F63EE41CF049D80F2B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"46AB5D56747C33F9052911BD";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"75DFFB9036C2D7F63EE41CF049D80F2B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 927 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"46AB5D56747C33F9052911BD") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F89A76077C769274434E7DE5C5C82829") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"46AB5D56747C33F9052911BD";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F89A76077C769274434E7DE5C5C82829") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 928 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"46AB5D56747C33F9052911BD") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2C7742EB276738CFE248879EE1D398B8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"46AB5D56747C33F9052911BD";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2C7742EB276738CFE248879EE1D398B8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 929 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"46AB5D56747C33F9052911BD") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BD3A5AD1EEFB39C205EDBFDE70A45457") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"46AB5D56747C33F9052911BD";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BD3A5AD1EEFB39C205EDBFDE70A45457") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 930 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"46AB5D56747C33F9052911BD") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9F88212393FE1E6753EB52D5898332B8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"46AB5D56747C33F9052911BD";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9F88212393FE1E6753EB52D5898332B8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 931 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"46AB5D56747C33F9052911BD") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0AF9DCCD4EE2D0C6F5F83B97B672A0FB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"46AB5D56747C33F9052911BD";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0AF9DCCD4EE2D0C6F5F83B97B672A0FB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 932 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"46AB5D56747C33F9052911BD") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BB69D0D588ADE17DAA0BC4BA5CD52FE3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"46AB5D56747C33F9052911BD";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BB69D0D588ADE17DAA0BC4BA5CD52FE3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 933 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"46AB5D56747C33F9052911BD") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"08611039E1E9FE9C6DEDA8B3481A8531") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"46AB5D56747C33F9052911BD";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"08611039E1E9FE9C6DEDA8B3481A8531") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 934 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"46AB5D56747C33F9052911BD") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D46D7BB1F9F6BFCB091A3FBFEAFD75A8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"46AB5D56747C33F9052911BD";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D46D7BB1F9F6BFCB091A3FBFEAFD75A8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 935 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"46AB5D56747C33F9052911BD") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6475A0EB2F51B68A4820F8BD7511EF93") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"46AB5D56747C33F9052911BD";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6475A0EB2F51B68A4820F8BD7511EF93") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 936 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"46AB5D56747C33F9052911BD") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1B7A49BFD31349A9C3B594351462C4F7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"46AB5D56747C33F9052911BD";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1B7A49BFD31349A9C3B594351462C4F7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 937 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"46AB5D56747C33F9052911BD") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"80BF81003159667CB1AF06CE96FC8F55") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"46AB5D56747C33F9052911BD";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"80BF81003159667CB1AF06CE96FC8F55") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 938 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"46AB5D56747C33F9052911BD") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EC07013486EFF692C19FA66282D4E6B0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"46AB5D56747C33F9052911BD";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EC07013486EFF692C19FA66282D4E6B0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 939 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"46AB5D56747C33F9052911BD") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B363AC4D9BCB8DA5E4F3CD2225BC9175") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"46AB5D56747C33F9052911BD";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B363AC4D9BCB8DA5E4F3CD2225BC9175") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 940 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"46AB5D56747C33F9052911BD") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F527DF4F87E927607E53FA8E4B9E1583") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"46AB5D56747C33F9052911BD";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F527DF4F87E927607E53FA8E4B9E1583") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 941 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"46AB5D56747C33F9052911BD") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5001E3B64EA9B4B4750634EDADBD2407") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"46AB5D56747C33F9052911BD";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5001E3B64EA9B4B4750634EDADBD2407") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 942 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"46AB5D56747C33F9052911BD") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4A7002B1942203618F7B75C72684DB3B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"46AB5D56747C33F9052911BD";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4A7002B1942203618F7B75C72684DB3B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 943 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"46AB5D56747C33F9052911BD") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3B919F060D1BAF52F78040C2D523ACBA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"46AB5D56747C33F9052911BD";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3B919F060D1BAF52F78040C2D523ACBA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 944 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"46AB5D56747C33F9052911BD") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F1DC1318A5B0D9B987346386D406DDCF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"46AB5D56747C33F9052911BD";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F1DC1318A5B0D9B987346386D406DDCF") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 945 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"46AB5D56747C33F9052911BD") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"795DE94B5C8ADB3A1F6797480FF2029E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"46AB5D56747C33F9052911BD";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"795DE94B5C8ADB3A1F6797480FF2029E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 946 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"46AB5D56747C33F9052911BD") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"65038953BA77306DC01D842A046BB46D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"46AB5D56747C33F9052911BD";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"65038953BA77306DC01D842A046BB46D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 947 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"46AB5D56747C33F9052911BD") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"94D5BBEFBC1DABB45AA1AC95897AB596") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"46AB5D56747C33F9052911BD";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"94D5BBEFBC1DABB45AA1AC95897AB596") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 948 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"46AB5D56747C33F9052911BD") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9BAB9C925761455519B93D21F58436B3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"46AB5D56747C33F9052911BD";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9BAB9C925761455519B93D21F58436B3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 949 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"46AB5D56747C33F9052911BD") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7D002DEECEC166BCC93DF940331DB4BD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"46AB5D56747C33F9052911BD";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7D002DEECEC166BCC93DF940331DB4BD") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 950 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"46AB5D56747C33F9052911BD") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BFA21E2D520B2924412C672B04C7FF8D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"46AB5D56747C33F9052911BD";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BFA21E2D520B2924412C672B04C7FF8D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 951 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"46AB5D56747C33F9052911BD") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1B6ECE03A8EF8FDDE730C35FD005CD0E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"46AB5D56747C33F9052911BD";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1B6ECE03A8EF8FDDE730C35FD005CD0E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 952 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"46AB5D56747C33F9052911BD") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F901FC1E73AE7CDDEDBF2F2C5218F458") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"46AB5D56747C33F9052911BD";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F901FC1E73AE7CDDEDBF2F2C5218F458") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 953 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"46AB5D56747C33F9052911BD") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8527A50853659CE4C32E4AF076E4CF6C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"46AB5D56747C33F9052911BD";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8527A50853659CE4C32E4AF076E4CF6C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 954 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"46AB5D56747C33F9052911BD") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"92A0E0EED8EB5F3C2774EE6641280E82") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"46AB5D56747C33F9052911BD";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"92A0E0EED8EB5F3C2774EE6641280E82") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 955 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"46AB5D56747C33F9052911BD") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6A8E2BB44C62F764443A6385D4C3BE10") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"46AB5D56747C33F9052911BD";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6A8E2BB44C62F764443A6385D4C3BE10") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 956 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"46AB5D56747C33F9052911BD") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3EBAA6D162A93BD7127B539ED368F77C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"46AB5D56747C33F9052911BD";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3EBAA6D162A93BD7127B539ED368F77C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 957 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"46AB5D56747C33F9052911BD") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D8D71C6F16C04677E5B5609D763712F1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"46AB5D56747C33F9052911BD";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-11)) = x"101112131415161718191A1B") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D8D71C6F16C04677E5B5609D763712F1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 958 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"46AB5D56747C33F9052911BDEC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"847203133E670C7D272226772962F66E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"46AB5D56747C33F9052911BDEC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"847203133E670C7D272226772962F66E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 959 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"46AB5D56747C33F9052911BDEC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"72FE83465A78D432C028ACAFFF25254D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"46AB5D56747C33F9052911BDEC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"72FE83465A78D432C028ACAFFF25254D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 960 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"46AB5D56747C33F9052911BDEC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FFBB0ED110CC91B0BD82CDBA7335024F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"46AB5D56747C33F9052911BDEC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FFBB0ED110CC91B0BD82CDBA7335024F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 961 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"46AB5D56747C33F9052911BDEC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2B563A3D4BDD3B0B1C8437C1572EB2DE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"46AB5D56747C33F9052911BDEC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2B563A3D4BDD3B0B1C8437C1572EB2DE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 962 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"46AB5D56747C33F9052911BDEC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BA1B220782413A06FB210F81C6597E31") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"46AB5D56747C33F9052911BDEC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BA1B220782413A06FB210F81C6597E31") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 963 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"46AB5D56747C33F9052911BDEC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"98A959F5FF441DA3AD27E28A3F7E18DE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"46AB5D56747C33F9052911BDEC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"98A959F5FF441DA3AD27E28A3F7E18DE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 964 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"46AB5D56747C33F9052911BDEC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0DD8A41B2258D3020B348BC8008F8A9D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"46AB5D56747C33F9052911BDEC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0DD8A41B2258D3020B348BC8008F8A9D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 965 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"46AB5D56747C33F9052911BDEC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BC48A803E417E2B954C774E5EA280585") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"46AB5D56747C33F9052911BDEC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BC48A803E417E2B954C774E5EA280585") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 966 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"46AB5D56747C33F9052911BDEC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0F4068EF8D53FD58932118ECFEE7AF57") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"46AB5D56747C33F9052911BDEC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0F4068EF8D53FD58932118ECFEE7AF57") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 967 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"46AB5D56747C33F9052911BDEC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D34C0367954CBC0FF7D68FE05C005FCE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"46AB5D56747C33F9052911BDEC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D34C0367954CBC0FF7D68FE05C005FCE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 968 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"46AB5D56747C33F9052911BDEC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6354D83D43EBB54EB6EC48E2C3ECC5F5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"46AB5D56747C33F9052911BDEC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6354D83D43EBB54EB6EC48E2C3ECC5F5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 969 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"46AB5D56747C33F9052911BDEC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1C5B3169BFA94A6D3D79246AA29FEE91") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"46AB5D56747C33F9052911BDEC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1C5B3169BFA94A6D3D79246AA29FEE91") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 970 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"46AB5D56747C33F9052911BDEC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"879EF9D65DE365B84F63B6912001A533") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"46AB5D56747C33F9052911BDEC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"879EF9D65DE365B84F63B6912001A533") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 971 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"46AB5D56747C33F9052911BDEC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EB2679E2EA55F5563F53163D3429CCD6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"46AB5D56747C33F9052911BDEC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EB2679E2EA55F5563F53163D3429CCD6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 972 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"46AB5D56747C33F9052911BDEC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B442D49BF7718E611A3F7D7D9341BB13") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"46AB5D56747C33F9052911BDEC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B442D49BF7718E611A3F7D7D9341BB13") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 973 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"46AB5D56747C33F9052911BDEC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F206A799EB5324A4809F4AD1FD633FE5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"46AB5D56747C33F9052911BDEC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F206A799EB5324A4809F4AD1FD633FE5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 974 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"46AB5D56747C33F9052911BDEC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"57209B602213B7708BCA84B21B400E61") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"46AB5D56747C33F9052911BDEC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"57209B602213B7708BCA84B21B400E61") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 975 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"46AB5D56747C33F9052911BDEC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4D517A67F89800A571B7C5989079F15D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"46AB5D56747C33F9052911BDEC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4D517A67F89800A571B7C5989079F15D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 976 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"46AB5D56747C33F9052911BDEC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3CB0E7D061A1AC96094CF09D63DE86DC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"46AB5D56747C33F9052911BDEC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3CB0E7D061A1AC96094CF09D63DE86DC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 977 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"46AB5D56747C33F9052911BDEC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F6FD6BCEC90ADA7D79F8D3D962FBF7A9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"46AB5D56747C33F9052911BDEC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F6FD6BCEC90ADA7D79F8D3D962FBF7A9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 978 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"46AB5D56747C33F9052911BDEC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7E7C919D3030D8FEE1AB2717B90F28F8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"46AB5D56747C33F9052911BDEC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7E7C919D3030D8FEE1AB2717B90F28F8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 979 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"46AB5D56747C33F9052911BDEC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6222F185D6CD33A93ED13475B2969E0B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"46AB5D56747C33F9052911BDEC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6222F185D6CD33A93ED13475B2969E0B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 980 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"46AB5D56747C33F9052911BDEC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"93F4C339D0A7A870A46D1CCA3F879FF0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"46AB5D56747C33F9052911BDEC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"93F4C339D0A7A870A46D1CCA3F879FF0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 981 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"46AB5D56747C33F9052911BDEC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9C8AE4443BDB4691E7758D7E43791CD5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"46AB5D56747C33F9052911BDEC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9C8AE4443BDB4691E7758D7E43791CD5") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 982 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"46AB5D56747C33F9052911BDEC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7A215538A27B657837F1491F85E09EDB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"46AB5D56747C33F9052911BDEC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7A215538A27B657837F1491F85E09EDB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 983 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"46AB5D56747C33F9052911BDEC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B88366FB3EB12AE0BFE0D774B23AD5EB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"46AB5D56747C33F9052911BDEC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B88366FB3EB12AE0BFE0D774B23AD5EB") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 984 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"46AB5D56747C33F9052911BDEC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1C4FB6D5C4558C1919FC730066F8E768") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"46AB5D56747C33F9052911BDEC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1C4FB6D5C4558C1919FC730066F8E768") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 985 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"46AB5D56747C33F9052911BDEC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FE2084C81F147F1913739F73E4E5DE3E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"46AB5D56747C33F9052911BDEC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FE2084C81F147F1913739F73E4E5DE3E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 986 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"46AB5D56747C33F9052911BDEC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8206DDDE3FDF9F203DE2FAAFC019E50A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"46AB5D56747C33F9052911BDEC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8206DDDE3FDF9F203DE2FAAFC019E50A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 987 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"46AB5D56747C33F9052911BDEC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"95819838B4515CF8D9B85E39F7D524E4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"46AB5D56747C33F9052911BDEC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"95819838B4515CF8D9B85E39F7D524E4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 988 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"46AB5D56747C33F9052911BDEC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6DAF536220D8F4A0BAF6D3DA623E9476") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"46AB5D56747C33F9052911BDEC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6DAF536220D8F4A0BAF6D3DA623E9476") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 989 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"46AB5D56747C33F9052911BDEC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"399BDE070E133813ECB7E3C16595DD1A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"46AB5D56747C33F9052911BDEC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"399BDE070E133813ECB7E3C16595DD1A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 990 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"46AB5D56747C33F9052911BDEC") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DFF664B97A7A45B31B79D0C2C0CA3897") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"46AB5D56747C33F9052911BDEC";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-12)) = x"101112131415161718191A1B1C") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DFF664B97A7A45B31B79D0C2C0CA3897") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 991 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"46AB5D56747C33F9052911BDEC7D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D50CA415F274D895DB9038B22ACEF597") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"46AB5D56747C33F9052911BDEC7D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D50CA415F274D895DB9038B22ACEF597") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 992 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"46AB5D56747C33F9052911BDEC7D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"23802440966B00DA3C9AB26AFC8926B4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"46AB5D56747C33F9052911BDEC7D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"23802440966B00DA3C9AB26AFC8926B4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 993 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"46AB5D56747C33F9052911BDEC7D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AEC5A9D7DCDF45584130D37F709901B6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"46AB5D56747C33F9052911BDEC7D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AEC5A9D7DCDF45584130D37F709901B6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 994 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"46AB5D56747C33F9052911BDEC7D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7A289D3B87CEEFE3E03629045482B127") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"46AB5D56747C33F9052911BDEC7D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7A289D3B87CEEFE3E03629045482B127") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 995 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"46AB5D56747C33F9052911BDEC7D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EB6585014E52EEEE07931144C5F57DC8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"46AB5D56747C33F9052911BDEC7D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EB6585014E52EEEE07931144C5F57DC8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 996 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"46AB5D56747C33F9052911BDEC7D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C9D7FEF33357C94B5195FC4F3CD21B27") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"46AB5D56747C33F9052911BDEC7D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C9D7FEF33357C94B5195FC4F3CD21B27") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 997 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"46AB5D56747C33F9052911BDEC7D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5CA6031DEE4B07EAF786950D03238964") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"46AB5D56747C33F9052911BDEC7D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5CA6031DEE4B07EAF786950D03238964") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 998 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"46AB5D56747C33F9052911BDEC7D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"ED360F0528043651A8756A20E984067C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"46AB5D56747C33F9052911BDEC7D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"ED360F0528043651A8756A20E984067C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 999 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"46AB5D56747C33F9052911BDEC7D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5E3ECFE9414029B06F930629FD4BACAE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"46AB5D56747C33F9052911BDEC7D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5E3ECFE9414029B06F930629FD4BACAE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1000 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"46AB5D56747C33F9052911BDEC7D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8232A461595F68E70B6491255FAC5C37") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"46AB5D56747C33F9052911BDEC7D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8232A461595F68E70B6491255FAC5C37") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1001 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"46AB5D56747C33F9052911BDEC7D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"322A7F3B8FF861A64A5E5627C040C60C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"46AB5D56747C33F9052911BDEC7D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"322A7F3B8FF861A64A5E5627C040C60C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1002 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"46AB5D56747C33F9052911BDEC7D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4D25966F73BA9E85C1CB3AAFA133ED68") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"46AB5D56747C33F9052911BDEC7D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4D25966F73BA9E85C1CB3AAFA133ED68") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1003 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"46AB5D56747C33F9052911BDEC7D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D6E05ED091F0B150B3D1A85423ADA6CA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"46AB5D56747C33F9052911BDEC7D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D6E05ED091F0B150B3D1A85423ADA6CA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1004 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"46AB5D56747C33F9052911BDEC7D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BA58DEE4264621BEC3E108F83785CF2F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"46AB5D56747C33F9052911BDEC7D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BA58DEE4264621BEC3E108F83785CF2F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1005 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"46AB5D56747C33F9052911BDEC7D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E53C739D3B625A89E68D63B890EDB8EA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"46AB5D56747C33F9052911BDEC7D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E53C739D3B625A89E68D63B890EDB8EA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1006 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"46AB5D56747C33F9052911BDEC7D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A378009F2740F04C7C2D5414FECF3C1C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"46AB5D56747C33F9052911BDEC7D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A378009F2740F04C7C2D5414FECF3C1C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1007 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"46AB5D56747C33F9052911BDEC7D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"065E3C66EE00639877789A7718EC0D98") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"46AB5D56747C33F9052911BDEC7D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"065E3C66EE00639877789A7718EC0D98") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1008 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"46AB5D56747C33F9052911BDEC7D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1C2FDD61348BD44D8D05DB5D93D5F2A4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"46AB5D56747C33F9052911BDEC7D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1C2FDD61348BD44D8D05DB5D93D5F2A4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1009 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"46AB5D56747C33F9052911BDEC7D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6DCE40D6ADB2787EF5FEEE5860728525") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"46AB5D56747C33F9052911BDEC7D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6DCE40D6ADB2787EF5FEEE5860728525") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1010 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"46AB5D56747C33F9052911BDEC7D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A783CCC805190E95854ACD1C6157F450") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"46AB5D56747C33F9052911BDEC7D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"A783CCC805190E95854ACD1C6157F450") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1011 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"46AB5D56747C33F9052911BDEC7D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2F02369BFC230C161D1939D2BAA32B01") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"46AB5D56747C33F9052911BDEC7D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2F02369BFC230C161D1939D2BAA32B01") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1012 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"46AB5D56747C33F9052911BDEC7D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"335C56831ADEE741C2632AB0B13A9DF2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"46AB5D56747C33F9052911BDEC7D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"335C56831ADEE741C2632AB0B13A9DF2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1013 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"46AB5D56747C33F9052911BDEC7D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C28A643F1CB47C9858DF020F3C2B9C09") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"46AB5D56747C33F9052911BDEC7D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C28A643F1CB47C9858DF020F3C2B9C09") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1014 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"46AB5D56747C33F9052911BDEC7D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CDF44342F7C892791BC793BB40D51F2C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"46AB5D56747C33F9052911BDEC7D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CDF44342F7C892791BC793BB40D51F2C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1015 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"46AB5D56747C33F9052911BDEC7D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2B5FF23E6E68B190CB4357DA864C9D22") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"46AB5D56747C33F9052911BDEC7D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2B5FF23E6E68B190CB4357DA864C9D22") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1016 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"46AB5D56747C33F9052911BDEC7D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E9FDC1FDF2A2FE084352C9B1B196D612") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"46AB5D56747C33F9052911BDEC7D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E9FDC1FDF2A2FE084352C9B1B196D612") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1017 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"46AB5D56747C33F9052911BDEC7D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4D3111D3084658F1E54E6DC56554E491") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"46AB5D56747C33F9052911BDEC7D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4D3111D3084658F1E54E6DC56554E491") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1018 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"46AB5D56747C33F9052911BDEC7D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AF5E23CED307ABF1EFC181B6E749DDC7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"46AB5D56747C33F9052911BDEC7D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AF5E23CED307ABF1EFC181B6E749DDC7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1019 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"46AB5D56747C33F9052911BDEC7D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D3787AD8F3CC4BC8C150E46AC3B5E6F3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"46AB5D56747C33F9052911BDEC7D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D3787AD8F3CC4BC8C150E46AC3B5E6F3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1020 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"46AB5D56747C33F9052911BDEC7D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C4FF3F3E78428810250A40FCF479271D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"46AB5D56747C33F9052911BDEC7D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"C4FF3F3E78428810250A40FCF479271D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1021 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"46AB5D56747C33F9052911BDEC7D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3CD1F464ECCB20484644CD1F6192978F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"46AB5D56747C33F9052911BDEC7D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3CD1F464ECCB20484644CD1F6192978F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1022 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"46AB5D56747C33F9052911BDEC7D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"68E57901C200ECFB1005FD046639DEE3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"46AB5D56747C33F9052911BDEC7D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"68E57901C200ECFB1005FD046639DEE3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1023 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"46AB5D56747C33F9052911BDEC7D") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8E88C3BFB669915BE7CBCE07C3663B6E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"46AB5D56747C33F9052911BDEC7D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-13)) = x"101112131415161718191A1B1C1D") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8E88C3BFB669915BE7CBCE07C3663B6E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1024 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"46AB5D56747C33F9052911BDEC7DB9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"84CBCA63C1F9391FF3CA70A5E9B8AC83") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"46AB5D56747C33F9052911BDEC7DB9";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"84CBCA63C1F9391FF3CA70A5E9B8AC83") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1025 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"46AB5D56747C33F9052911BDEC7DB9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"72474A36A5E6E15014C0FA7D3FFF7FA0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"46AB5D56747C33F9052911BDEC7DB9";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"72474A36A5E6E15014C0FA7D3FFF7FA0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1026 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"46AB5D56747C33F9052911BDEC7DB9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FF02C7A1EF52A4D2696A9B68B3EF58A2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"46AB5D56747C33F9052911BDEC7DB9";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FF02C7A1EF52A4D2696A9B68B3EF58A2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1027 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"46AB5D56747C33F9052911BDEC7DB9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2BEFF34DB4430E69C86C611397F4E833") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"46AB5D56747C33F9052911BDEC7DB9";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"2BEFF34DB4430E69C86C611397F4E833") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1028 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"46AB5D56747C33F9052911BDEC7DB9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BAA2EB777DDF0F642FC95953068324DC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"46AB5D56747C33F9052911BDEC7DB9";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BAA2EB777DDF0F642FC95953068324DC") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1029 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"46AB5D56747C33F9052911BDEC7DB9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9810908500DA28C179CFB458FFA44233") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"46AB5D56747C33F9052911BDEC7DB9";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9810908500DA28C179CFB458FFA44233") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1030 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"46AB5D56747C33F9052911BDEC7DB9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0D616D6BDDC6E660DFDCDD1AC055D070") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"46AB5D56747C33F9052911BDEC7DB9";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0D616D6BDDC6E660DFDCDD1AC055D070") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1031 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"46AB5D56747C33F9052911BDEC7DB9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BCF161731B89D7DB802F22372AF25F68") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"46AB5D56747C33F9052911BDEC7DB9";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"BCF161731B89D7DB802F22372AF25F68") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1032 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"46AB5D56747C33F9052911BDEC7DB9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0FF9A19F72CDC83A47C94E3E3E3DF5BA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"46AB5D56747C33F9052911BDEC7DB9";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0FF9A19F72CDC83A47C94E3E3E3DF5BA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1033 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"46AB5D56747C33F9052911BDEC7DB9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D3F5CA176AD2896D233ED9329CDA0523") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"46AB5D56747C33F9052911BDEC7DB9";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"D3F5CA176AD2896D233ED9329CDA0523") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1034 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"46AB5D56747C33F9052911BDEC7DB9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"63ED114DBC75802C62041E3003369F18") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"46AB5D56747C33F9052911BDEC7DB9";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"63ED114DBC75802C62041E3003369F18") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1035 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"46AB5D56747C33F9052911BDEC7DB9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1CE2F81940377F0FE99172B86245B47C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"46AB5D56747C33F9052911BDEC7DB9";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1CE2F81940377F0FE99172B86245B47C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1036 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"46AB5D56747C33F9052911BDEC7DB9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"872730A6A27D50DA9B8BE043E0DBFFDE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"46AB5D56747C33F9052911BDEC7DB9";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"872730A6A27D50DA9B8BE043E0DBFFDE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1037 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"46AB5D56747C33F9052911BDEC7DB9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EB9FB09215CBC034EBBB40EFF4F3963B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"46AB5D56747C33F9052911BDEC7DB9";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EB9FB09215CBC034EBBB40EFF4F3963B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1038 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"46AB5D56747C33F9052911BDEC7DB9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B4FB1DEB08EFBB03CED72BAF539BE1FE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"46AB5D56747C33F9052911BDEC7DB9";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B4FB1DEB08EFBB03CED72BAF539BE1FE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1039 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"46AB5D56747C33F9052911BDEC7DB9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F2BF6EE914CD11C654771C033DB96508") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"46AB5D56747C33F9052911BDEC7DB9";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F2BF6EE914CD11C654771C033DB96508") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1040 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"46AB5D56747C33F9052911BDEC7DB9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"57995210DD8D82125F22D260DB9A548C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"46AB5D56747C33F9052911BDEC7DB9";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"57995210DD8D82125F22D260DB9A548C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1041 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"46AB5D56747C33F9052911BDEC7DB9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4DE8B317070635C7A55F934A50A3ABB0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"46AB5D56747C33F9052911BDEC7DB9";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"4DE8B317070635C7A55F934A50A3ABB0") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1042 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"46AB5D56747C33F9052911BDEC7DB9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3C092EA09E3F99F4DDA4A64FA304DC31") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"46AB5D56747C33F9052911BDEC7DB9";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"3C092EA09E3F99F4DDA4A64FA304DC31") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1043 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"46AB5D56747C33F9052911BDEC7DB9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F644A2BE3694EF1FAD10850BA221AD44") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"46AB5D56747C33F9052911BDEC7DB9";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"F644A2BE3694EF1FAD10850BA221AD44") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1044 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"46AB5D56747C33F9052911BDEC7DB9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7EC558EDCFAEED9C354371C579D57215") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"46AB5D56747C33F9052911BDEC7DB9";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7EC558EDCFAEED9C354371C579D57215") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1045 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"46AB5D56747C33F9052911BDEC7DB9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"629B38F5295306CBEA3962A7724CC4E6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"46AB5D56747C33F9052911BDEC7DB9";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"629B38F5295306CBEA3962A7724CC4E6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1046 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"46AB5D56747C33F9052911BDEC7DB9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"934D0A492F399D1270854A18FF5DC51D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"46AB5D56747C33F9052911BDEC7DB9";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"934D0A492F399D1270854A18FF5DC51D") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1047 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"46AB5D56747C33F9052911BDEC7DB9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9C332D34C44573F3339DDBAC83A34638") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"46AB5D56747C33F9052911BDEC7DB9";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9C332D34C44573F3339DDBAC83A34638") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1048 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"46AB5D56747C33F9052911BDEC7DB9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7A989C485DE5501AE3191FCD453AC436") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"46AB5D56747C33F9052911BDEC7DB9";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7A989C485DE5501AE3191FCD453AC436") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1049 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"46AB5D56747C33F9052911BDEC7DB9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B83AAF8BC12F1F826B0881A672E08F06") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"46AB5D56747C33F9052911BDEC7DB9";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B83AAF8BC12F1F826B0881A672E08F06") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1050 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"46AB5D56747C33F9052911BDEC7DB9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1CF67FA53BCBB97BCD1425D2A622BD85") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"46AB5D56747C33F9052911BDEC7DB9";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1CF67FA53BCBB97BCD1425D2A622BD85") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1051 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"46AB5D56747C33F9052911BDEC7DB9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FE994DB8E08A4A7BC79BC9A1243F84D3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"46AB5D56747C33F9052911BDEC7DB9";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FE994DB8E08A4A7BC79BC9A1243F84D3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1052 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"46AB5D56747C33F9052911BDEC7DB9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"82BF14AEC041AA42E90AAC7D00C3BFE7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"46AB5D56747C33F9052911BDEC7DB9";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"82BF14AEC041AA42E90AAC7D00C3BFE7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1053 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"46AB5D56747C33F9052911BDEC7DB9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"953851484BCF699A0D5008EB370F7E09") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"46AB5D56747C33F9052911BDEC7DB9";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"953851484BCF699A0D5008EB370F7E09") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1054 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"46AB5D56747C33F9052911BDEC7DB9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6D169A12DF46C1C26E1E8508A2E4CE9B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"46AB5D56747C33F9052911BDEC7DB9";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6D169A12DF46C1C26E1E8508A2E4CE9B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1055 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"46AB5D56747C33F9052911BDEC7DB9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"39221777F18D0D71385FB513A54F87F7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"46AB5D56747C33F9052911BDEC7DB9";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"39221777F18D0D71385FB513A54F87F7") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1056 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"46AB5D56747C33F9052911BDEC7DB9") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DF4FADC985E470D1CF9186100010627A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"46AB5D56747C33F9052911BDEC7DB9";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-14)) = x"101112131415161718191A1B1C1D1E") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DF4FADC985E470D1CF9186100010627A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1057 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"A04A9135204535AE92BD5D11629F3C8F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"63C450C2B5ED4EAABDD2360D20946B01") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"A04A9135204535AE92BD5D11629F3C8F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"63C450C2B5ED4EAABDD2360D20946B01") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1058 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"A04A9135204535AE92BD5D11629F3C8F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9548D097D1F296E55AD8BCD5F6D3B822") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"00";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"A04A9135204535AE92BD5D11629F3C8F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9548D097D1F296E55AD8BCD5F6D3B822") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1059 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"A04A9135204535AE92BD5D11629F3C8F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"180D5D009B46D3672772DDC07AC39F20") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"0001";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"A04A9135204535AE92BD5D11629F3C8F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"180D5D009B46D3672772DDC07AC39F20") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1060 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"A04A9135204535AE92BD5D11629F3C8F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CCE069ECC05779DC867427BB5ED82FB1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"000102";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"A04A9135204535AE92BD5D11629F3C8F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"CCE069ECC05779DC867427BB5ED82FB1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1061 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"A04A9135204535AE92BD5D11629F3C8F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5DAD71D609CB78D161D11FFBCFAFE35E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"00010203";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"A04A9135204535AE92BD5D11629F3C8F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5DAD71D609CB78D161D11FFBCFAFE35E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1062 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"A04A9135204535AE92BD5D11629F3C8F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7F1F0A2474CE5F7437D7F2F0368885B1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"0001020304";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"A04A9135204535AE92BD5D11629F3C8F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7F1F0A2474CE5F7437D7F2F0368885B1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1063 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"A04A9135204535AE92BD5D11629F3C8F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EA6EF7CAA9D291D591C49BB2097917F2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"000102030405";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"A04A9135204535AE92BD5D11629F3C8F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"EA6EF7CAA9D291D591C49BB2097917F2") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1064 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"A04A9135204535AE92BD5D11629F3C8F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5BFEFBD26F9DA06ECE37649FE3DE98EA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"00010203040506";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"A04A9135204535AE92BD5D11629F3C8F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5BFEFBD26F9DA06ECE37649FE3DE98EA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1065 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"A04A9135204535AE92BD5D11629F3C8F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E8F63B3E06D9BF8F09D10896F7113238") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"0001020304050607";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"A04A9135204535AE92BD5D11629F3C8F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"E8F63B3E06D9BF8F09D10896F7113238") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1066 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"A04A9135204535AE92BD5D11629F3C8F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"34FA50B61EC6FED86D269F9A55F6C2A1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"000102030405060708";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"A04A9135204535AE92BD5D11629F3C8F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"34FA50B61EC6FED86D269F9A55F6C2A1") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1067 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"A04A9135204535AE92BD5D11629F3C8F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"84E28BECC861F7992C1C5898CA1A589A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"00010203040506070809";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"A04A9135204535AE92BD5D11629F3C8F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"84E28BECC861F7992C1C5898CA1A589A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1068 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"A04A9135204535AE92BD5D11629F3C8F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FBED62B8342308BAA7893410AB6973FE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"000102030405060708090A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"A04A9135204535AE92BD5D11629F3C8F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FBED62B8342308BAA7893410AB6973FE") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1069 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"A04A9135204535AE92BD5D11629F3C8F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6028AA07D669276FD593A6EB29F7385C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"000102030405060708090A0B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"A04A9135204535AE92BD5D11629F3C8F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"6028AA07D669276FD593A6EB29F7385C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1070 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"A04A9135204535AE92BD5D11629F3C8F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0C902A3361DFB781A5A306473DDF51B9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"000102030405060708090A0B0C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"A04A9135204535AE92BD5D11629F3C8F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"0C902A3361DFB781A5A306473DDF51B9") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1071 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"A04A9135204535AE92BD5D11629F3C8F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"53F4874A7CFBCCB680CF6D079AB7267C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"000102030405060708090A0B0C0D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"A04A9135204535AE92BD5D11629F3C8F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"53F4874A7CFBCCB680CF6D079AB7267C") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1072 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"A04A9135204535AE92BD5D11629F3C8F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"15B0F44860D966731A6F5AABF495A28A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"000102030405060708090A0B0C0D0E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"A04A9135204535AE92BD5D11629F3C8F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"15B0F44860D966731A6F5AABF495A28A") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1073 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"A04A9135204535AE92BD5D11629F3C8F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B096C8B1A999F5A7113A94C812B6930E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"A04A9135204535AE92BD5D11629F3C8F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"B096C8B1A999F5A7113A94C812B6930E") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1074 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"A04A9135204535AE92BD5D11629F3C8F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AAE729B673124272EB47D5E2998F6C32") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-0)) <= x"10";
      Block_Size <= x"0";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"A04A9135204535AE92BD5D11629F3C8F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"AAE729B673124272EB47D5E2998F6C32") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1075 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"A04A9135204535AE92BD5D11629F3C8F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DB06B401EA2BEE4193BCE0E76A281BB3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-1)) <= x"1011";
      Block_Size <= x"1";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"A04A9135204535AE92BD5D11629F3C8F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DB06B401EA2BEE4193BCE0E76A281BB3") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1076 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"A04A9135204535AE92BD5D11629F3C8F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"114B381F428098AAE308C3A36B0D6AC6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-2)) <= x"101112";
      Block_Size <= x"2";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"A04A9135204535AE92BD5D11629F3C8F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"114B381F428098AAE308C3A36B0D6AC6") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1077 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"A04A9135204535AE92BD5D11629F3C8F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"99CAC24CBBBA9A297B5B376DB0F9B597") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-3)) <= x"10111213";
      Block_Size <= x"3";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"A04A9135204535AE92BD5D11629F3C8F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"99CAC24CBBBA9A297B5B376DB0F9B597") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1078 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"A04A9135204535AE92BD5D11629F3C8F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8594A2545D47717EA421240FBB600364") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-4)) <= x"1011121314";
      Block_Size <= x"4";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"A04A9135204535AE92BD5D11629F3C8F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8594A2545D47717EA421240FBB600364") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1079 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"A04A9135204535AE92BD5D11629F3C8F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"744290E85B2DEAA73E9D0CB03671029F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-5)) <= x"101112131415";
      Block_Size <= x"5";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"A04A9135204535AE92BD5D11629F3C8F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"744290E85B2DEAA73E9D0CB03671029F") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1080 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"A04A9135204535AE92BD5D11629F3C8F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7B3CB795B05104467D859D044A8F81BA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-6)) <= x"10111213141516";
      Block_Size <= x"6";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"A04A9135204535AE92BD5D11629F3C8F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7B3CB795B05104467D859D044A8F81BA") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1081 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"A04A9135204535AE92BD5D11629F3C8F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9D9706E929F127AFAD0159658C1603B4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-7)) <= x"1011121314151617";
      Block_Size <= x"7";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"A04A9135204535AE92BD5D11629F3C8F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"9D9706E929F127AFAD0159658C1603B4") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1082 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"A04A9135204535AE92BD5D11629F3C8F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5F35352AB53B68372510C70EBBCC4884") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-8)) <= x"101112131415161718";
      Block_Size <= x"8";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"A04A9135204535AE92BD5D11629F3C8F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"5F35352AB53B68372510C70EBBCC4884") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1083 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"A04A9135204535AE92BD5D11629F3C8F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FBF9E5044FDFCECE830C637A6F0E7A07") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-9)) <= x"10111213141516171819";
      Block_Size <= x"9";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"A04A9135204535AE92BD5D11629F3C8F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"FBF9E5044FDFCECE830C637A6F0E7A07") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1084 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"A04A9135204535AE92BD5D11629F3C8F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1996D719949E3DCE89838F09ED134351") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-10)) <= x"101112131415161718191A";
      Block_Size <= x"a";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"A04A9135204535AE92BD5D11629F3C8F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"1996D719949E3DCE89838F09ED134351") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1085 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"A04A9135204535AE92BD5D11629F3C8F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"65B08E0FB455DDF7A712EAD5C9EF7865") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-11)) <= x"101112131415161718191A1B";
      Block_Size <= x"b";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"A04A9135204535AE92BD5D11629F3C8F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"65B08E0FB455DDF7A712EAD5C9EF7865") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1086 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"A04A9135204535AE92BD5D11629F3C8F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7237CBE93FDB1E2F43484E43FE23B98B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-12)) <= x"101112131415161718191A1B1C";
      Block_Size <= x"c";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"A04A9135204535AE92BD5D11629F3C8F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"7237CBE93FDB1E2F43484E43FE23B98B") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1087 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"A04A9135204535AE92BD5D11629F3C8F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8A1900B3AB52B6772006C3A06BC80919") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-13)) <= x"101112131415161718191A1B1C1D";
      Block_Size <= x"d";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"A04A9135204535AE92BD5D11629F3C8F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"8A1900B3AB52B6772006C3A06BC80919") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1088 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"A04A9135204535AE92BD5D11629F3C8F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DE2D8DD685997AC47647F3BB6C634075") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-14)) <= x"101112131415161718191A1B1C1D1E";
      Block_Size <= x"e";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"A04A9135204535AE92BD5D11629F3C8F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"DE2D8DD685997AC47647F3BB6C634075") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      --------- test no. 1089 ----------

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"141DE4122F09D2E045E60CF3C96B1534") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      enc <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"A04A9135204535AE92BD5D11629F3C8F") then
         report "---- Encryption Passed -----";
      else
         report "**** Encryption Failed *****";
      end if;

      wait for clk_period * 1;
      enc <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"38403768F1F007648189C0B8C93CA5F8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --=======================================================================================

      rst     <= '1';
      a_data  <= '0';
      enc     <= '0';
      dec     <= '0';
      gen_tag <= '0';
      K       <= x"000102030405060708090A0B0C0D0E0F";
      N       <= x"000102030405060708090A0B";
      wait for clk_period * 1;

      rst <= '0';
      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"000102030405060708090A0B0C0D0E0F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      a_data <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"101112131415161718191A1B1C1D1E1F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      wait for clk_period * 1;
      a_data <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"141DE4122F09D2E045E60CF3C96B1534";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"000102030405060708090A0B0C0D0E0F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      dec <= '1';
      Input(8*16-1 downto 8*(15-15)) <= x"A04A9135204535AE92BD5D11629F3C8F";
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Output(8*16-1 downto 8*(15-15)) = x"101112131415161718191A1B1C1D1E1F") then
         report "---- Decryption Passed -----";
      else
         report "**** Decryption Failed *****";
      end if;

      wait for clk_period * 1;
      dec <= '0';
      wait for clk_period * 1;

      gen_tag <= '1';
      Block_Size <= x"f";

      wait until done = '1';
      wait for clk_period*0.5;

      if (Tag = x"38403768F1F007648189C0B8C93CA5F8") then
      	 report "------------ Tag Passed -----";
      else
      	 report "************ Tag Failed *****";
      end if;

      --======================================================================================= 

      wait;
   end process;

END;
